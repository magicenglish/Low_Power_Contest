
module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   N23, ld_r, N34, N35, N36, N37, N38, N39, N40, N41, N50, N51, N52, N53,
         N54, N55, N56, N57, N66, N67, N68, N69, N70, N71, N72, N73, N82, N83,
         N84, N85, N86, N87, N88, N89, N98, N99, N100, N101, N102, N103, N104,
         N105, N114, N115, N116, N117, N118, N119, N120, N121, N130, N131,
         N132, N133, N134, N135, N136, N137, N146, N147, N148, N149, N150,
         N151, N152, N153, N162, N163, N164, N165, N166, N167, N168, N169,
         N178, N179, N180, N181, N182, N183, N184, N185, N194, N195, N196,
         N197, N198, N199, N200, N201, N210, N211, N212, N213, N214, N215,
         N216, N217, N226, N227, N228, N229, N230, N231, N232, N233, N242,
         N243, N244, N245, N246, N247, N248, N249, N258, N259, N260, N261,
         N262, N263, N264, N265, N274, N275, N276, N277, N278, N279, N280,
         N281, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, \u0/N271 , \u0/N270 ,
         \u0/N269 , \u0/N268 , \u0/N267 , \u0/N266 , \u0/N265 , \u0/N264 ,
         \u0/N263 , \u0/N262 , \u0/N261 , \u0/N260 , \u0/N259 , \u0/N258 ,
         \u0/N257 , \u0/N256 , \u0/N255 , \u0/N254 , \u0/N253 , \u0/N252 ,
         \u0/N251 , \u0/N250 , \u0/N249 , \u0/N248 , \u0/N247 , \u0/N246 ,
         \u0/N245 , \u0/N244 , \u0/N243 , \u0/N242 , \u0/N241 , \u0/N240 ,
         \u0/N205 , \u0/N204 , \u0/N203 , \u0/N202 , \u0/N201 , \u0/N200 ,
         \u0/N199 , \u0/N198 , \u0/N197 , \u0/N196 , \u0/N195 , \u0/N194 ,
         \u0/N193 , \u0/N192 , \u0/N191 , \u0/N190 , \u0/N189 , \u0/N188 ,
         \u0/N187 , \u0/N186 , \u0/N185 , \u0/N184 , \u0/N183 , \u0/N182 ,
         \u0/N181 , \u0/N180 , \u0/N179 , \u0/N178 , \u0/N177 , \u0/N176 ,
         \u0/N175 , \u0/N174 , \u0/N139 , \u0/N138 , \u0/N137 , \u0/N136 ,
         \u0/N135 , \u0/N134 , \u0/N133 , \u0/N132 , \u0/N131 , \u0/N130 ,
         \u0/N129 , \u0/N128 , \u0/N127 , \u0/N126 , \u0/N125 , \u0/N124 ,
         \u0/N123 , \u0/N122 , \u0/N121 , \u0/N120 , \u0/N119 , \u0/N118 ,
         \u0/N117 , \u0/N116 , \u0/N115 , \u0/N114 , \u0/N113 , \u0/N112 ,
         \u0/N111 , \u0/N110 , \u0/N109 , \u0/N108 , \u0/N73 , \u0/N72 ,
         \u0/N71 , \u0/N70 , \u0/N69 , \u0/N68 , \u0/N67 , \u0/N66 , \u0/N65 ,
         \u0/N64 , \u0/N63 , \u0/N62 , \u0/N61 , \u0/N60 , \u0/N59 , \u0/N58 ,
         \u0/N57 , \u0/N56 , \u0/N55 , \u0/N54 , \u0/N53 , \u0/N52 , \u0/N51 ,
         \u0/N50 , \u0/N49 , \u0/N48 , \u0/N47 , \u0/N46 , \u0/N45 , \u0/N44 ,
         \u0/N43 , \u0/N42 , \u0/r0/N81 , \u0/r0/N80 , \u0/r0/N79 ,
         \u0/r0/N78 , \u0/r0/N77 , \u0/r0/N76 , \u0/r0/N75 , \u0/r0/N74 ,
         \u0/r0/N73 , \u0/r0/N72 , \u0/r0/N71 , \u0/r0/N70 , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n7664, n7665, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa23;
  wire   [7:0] sa13;
  wire   [7:0] sa03;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa22;
  wire   [7:0] sa12;
  wire   [7:0] sa02;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa21;
  wire   [7:0] sa11;
  wire   [7:0] sa01;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa20;
  wire   [7:0] sa10;
  wire   [7:0] sa00;
  wire   [31:0] \u0/rcon ;
  wire   [3:0] \u0/r0/rcnt ;

  HS65_LL_DFPQX4 \sa30_reg[0]  ( .D(N226), .CP(clk), .Q(sa30[0]) );
  HS65_LL_DFPQX4 \sa33_reg[0]  ( .D(N34), .CP(clk), .Q(sa33[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][0]  ( .D(\u0/N174 ), .CP(clk), .Q(w2[0]) );
  HS65_LL_DFPQX4 \sa32_reg[0]  ( .D(N98), .CP(clk), .Q(sa32[0]) );
  HS65_LL_DFPQX4 \sa31_reg[0]  ( .D(N162), .CP(clk), .Q(sa31[0]) );
  HS65_LL_DFPQX4 \sa30_reg[1]  ( .D(N227), .CP(clk), .Q(sa30[1]) );
  HS65_LL_DFPQX4 \sa33_reg[1]  ( .D(N35), .CP(clk), .Q(sa33[1]) );
  HS65_LL_DFPQX4 \sa30_reg[2]  ( .D(N228), .CP(clk), .Q(sa30[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][2]  ( .D(\u0/N242 ), .CP(clk), .Q(w3[2]) );
  HS65_LL_DFPQX4 \sa31_reg[2]  ( .D(N164), .CP(clk), .Q(sa31[2]) );
  HS65_LL_DFPQX4 \sa33_reg[3]  ( .D(N37), .CP(clk), .Q(sa33[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][3]  ( .D(\u0/N177 ), .CP(clk), .Q(w2[3]) );
  HS65_LL_DFPQX4 \sa32_reg[3]  ( .D(N101), .CP(clk), .Q(sa32[3]) );
  HS65_LL_DFPQX4 \sa31_reg[3]  ( .D(N165), .CP(clk), .Q(sa31[3]) );
  HS65_LL_DFPQX4 \sa30_reg[4]  ( .D(N230), .CP(clk), .Q(sa30[4]) );
  HS65_LL_DFPQX4 \sa33_reg[4]  ( .D(N38), .CP(clk), .Q(sa33[4]) );
  HS65_LL_DFPQX4 \sa32_reg[4]  ( .D(N102), .CP(clk), .Q(sa32[4]) );
  HS65_LL_DFPQX4 \sa31_reg[4]  ( .D(N166), .CP(clk), .Q(sa31[4]) );
  HS65_LL_DFPQX4 \sa33_reg[5]  ( .D(N39), .CP(clk), .Q(sa33[5]) );
  HS65_LL_DFPQX4 \sa32_reg[5]  ( .D(N103), .CP(clk), .Q(sa32[5]) );
  HS65_LL_DFPQX4 \sa30_reg[6]  ( .D(N232), .CP(clk), .Q(sa30[6]) );
  HS65_LL_DFPQX4 \sa33_reg[6]  ( .D(N40), .CP(clk), .Q(sa33[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][6]  ( .D(\u0/N180 ), .CP(clk), .Q(w2[6]) );
  HS65_LL_DFPQX4 \sa32_reg[6]  ( .D(N104), .CP(clk), .Q(sa32[6]) );
  HS65_LL_DFPQX4 \sa30_reg[7]  ( .D(N233), .CP(clk), .Q(sa30[7]) );
  HS65_LL_DFPQX4 \sa32_reg[7]  ( .D(N105), .CP(clk), .Q(sa32[7]) );
  HS65_LL_DFPQX4 \sa31_reg[7]  ( .D(N169), .CP(clk), .Q(sa31[7]) );
  HS65_LL_DFPQX4 \sa23_reg[0]  ( .D(N50), .CP(clk), .Q(sa23[0]) );
  HS65_LL_DFPQX4 \sa22_reg[0]  ( .D(N114), .CP(clk), .Q(sa22[0]) );
  HS65_LL_DFPQX4 \sa21_reg[0]  ( .D(N178), .CP(clk), .Q(sa21[0]) );
  HS65_LL_DFPQX4 \sa20_reg[1]  ( .D(N243), .CP(clk), .Q(sa20[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][9]  ( .D(\u0/N183 ), .CP(clk), .Q(w2[9]) );
  HS65_LL_DFPQX4 \sa22_reg[1]  ( .D(N115), .CP(clk), .Q(sa22[1]) );
  HS65_LL_DFPQX4 \sa20_reg[2]  ( .D(N244), .CP(clk), .Q(sa20[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][10]  ( .D(\u0/N184 ), .CP(clk), .Q(w2[10]) );
  HS65_LL_DFPQX4 \sa22_reg[2]  ( .D(N116), .CP(clk), .Q(sa22[2]) );
  HS65_LL_DFPQX4 \sa20_reg[3]  ( .D(N245), .CP(clk), .Q(sa20[3]) );
  HS65_LL_DFPQX4 \sa23_reg[3]  ( .D(N53), .CP(clk), .Q(sa23[3]) );
  HS65_LL_DFPQX4 \sa22_reg[3]  ( .D(N117), .CP(clk), .Q(sa22[3]) );
  HS65_LL_DFPQX4 \sa20_reg[4]  ( .D(N246), .CP(clk), .Q(sa20[4]) );
  HS65_LL_DFPQX4 \sa23_reg[4]  ( .D(N54), .CP(clk), .Q(sa23[4]) );
  HS65_LL_DFPQX4 \sa22_reg[4]  ( .D(N118), .CP(clk), .Q(sa22[4]) );
  HS65_LL_DFPQX4 \sa21_reg[4]  ( .D(N182), .CP(clk), .Q(sa21[4]) );
  HS65_LL_DFPQX4 \sa22_reg[5]  ( .D(N119), .CP(clk), .Q(sa22[5]) );
  HS65_LL_DFPQX4 \sa23_reg[6]  ( .D(N56), .CP(clk), .Q(sa23[6]) );
  HS65_LL_DFPQX4 \sa22_reg[6]  ( .D(N120), .CP(clk), .Q(sa22[6]) );
  HS65_LL_DFPQX4 \sa22_reg[7]  ( .D(N121), .CP(clk), .Q(sa22[7]) );
  HS65_LL_DFPQX4 \sa10_reg[0]  ( .D(N258), .CP(clk), .Q(sa10[0]) );
  HS65_LL_DFPQX4 \sa13_reg[0]  ( .D(N66), .CP(clk), .Q(sa13[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][16]  ( .D(\u0/N190 ), .CP(clk), .Q(w2[16]) );
  HS65_LL_DFPQX4 \sa12_reg[0]  ( .D(N130), .CP(clk), .Q(sa12[0]) );
  HS65_LL_DFPQX4 \sa11_reg[0]  ( .D(N194), .CP(clk), .Q(sa11[0]) );
  HS65_LL_DFPQX4 \sa10_reg[1]  ( .D(N259), .CP(clk), .Q(sa10[1]) );
  HS65_LL_DFPQX4 \sa13_reg[1]  ( .D(N67), .CP(clk), .Q(sa13[1]) );
  HS65_LL_DFPQX4 \sa10_reg[2]  ( .D(N260), .CP(clk), .Q(sa10[2]) );
  HS65_LL_DFPQX4 \sa13_reg[2]  ( .D(N68), .CP(clk), .Q(sa13[2]) );
  HS65_LL_DFPQX4 \sa12_reg[2]  ( .D(N132), .CP(clk), .Q(sa12[2]) );
  HS65_LL_DFPQX4 \sa11_reg[2]  ( .D(N196), .CP(clk), .Q(sa11[2]) );
  HS65_LL_DFPQX4 \sa10_reg[3]  ( .D(N261), .CP(clk), .Q(sa10[3]) );
  HS65_LL_DFPQX4 \sa13_reg[3]  ( .D(N69), .CP(clk), .Q(sa13[3]) );
  HS65_LL_DFPQX4 \sa12_reg[3]  ( .D(N133), .CP(clk), .Q(sa12[3]) );
  HS65_LL_DFPQX4 \sa11_reg[3]  ( .D(N197), .CP(clk), .Q(sa11[3]) );
  HS65_LL_DFPQX4 \sa10_reg[4]  ( .D(N262), .CP(clk), .Q(sa10[4]) );
  HS65_LL_DFPQX4 \sa13_reg[4]  ( .D(N70), .CP(clk), .Q(sa13[4]) );
  HS65_LL_DFPQX4 \sa12_reg[4]  ( .D(N134), .CP(clk), .Q(sa12[4]) );
  HS65_LL_DFPQX4 \sa11_reg[4]  ( .D(N198), .CP(clk), .Q(sa11[4]) );
  HS65_LL_DFPQX4 \sa13_reg[5]  ( .D(N71), .CP(clk), .Q(sa13[5]) );
  HS65_LL_DFPQX4 \sa11_reg[7]  ( .D(N201), .CP(clk), .Q(sa11[7]) );
  HS65_LL_DFPQX4 \sa03_reg[0]  ( .D(N82), .CP(clk), .Q(sa03[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][24]  ( .D(\u0/N198 ), .CP(clk), .Q(w2[24]) );
  HS65_LL_DFPQX4 \sa02_reg[0]  ( .D(N146), .CP(clk), .Q(sa02[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][24]  ( .D(\u0/N132 ), .CP(clk), .Q(w1[24]) );
  HS65_LL_DFPQX4 \sa01_reg[0]  ( .D(N210), .CP(clk), .Q(sa01[0]) );
  HS65_LL_DFPQX4 \sa00_reg[0]  ( .D(N274), .CP(clk), .Q(sa00[0]) );
  HS65_LL_DFPQX4 \sa03_reg[2]  ( .D(N84), .CP(clk), .Q(sa03[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][26]  ( .D(\u0/N200 ), .CP(clk), .Q(w2[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][26]  ( .D(\u0/N134 ), .CP(clk), .Q(w1[26]) );
  HS65_LL_DFPQX4 \sa01_reg[2]  ( .D(N212), .CP(clk), .Q(sa01[2]) );
  HS65_LL_DFPQX4 \sa00_reg[2]  ( .D(N276), .CP(clk), .Q(sa00[2]) );
  HS65_LL_DFPQX4 \sa03_reg[3]  ( .D(N85), .CP(clk), .Q(sa03[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][27]  ( .D(\u0/N201 ), .CP(clk), .Q(w2[27]) );
  HS65_LL_DFPQX4 \sa02_reg[3]  ( .D(N149), .CP(clk), .Q(sa02[3]) );
  HS65_LL_DFPQX4 \sa01_reg[3]  ( .D(N213), .CP(clk), .Q(sa01[3]) );
  HS65_LL_DFPQX4 \sa00_reg[3]  ( .D(N277), .CP(clk), .Q(sa00[3]) );
  HS65_LL_DFPQX4 \sa03_reg[4]  ( .D(N86), .CP(clk), .Q(sa03[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][28]  ( .D(\u0/N202 ), .CP(clk), .Q(w2[28]) );
  HS65_LL_DFPQX4 \sa02_reg[4]  ( .D(N150), .CP(clk), .Q(sa02[4]) );
  HS65_LL_DFPQX4 \sa01_reg[4]  ( .D(N214), .CP(clk), .Q(sa01[4]) );
  HS65_LL_DFPQX4 \sa00_reg[4]  ( .D(N278), .CP(clk), .Q(sa00[4]) );
  HS65_LL_DFPQX4 \sa00_reg[5]  ( .D(N279), .CP(clk), .Q(sa00[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][30]  ( .D(\u0/N204 ), .CP(clk), .Q(w2[30]) );
  HS65_LL_DFPQX4 \sa00_reg[6]  ( .D(N280), .CP(clk), .Q(sa00[6]) );
  HS65_LL_DFPQX4 \sa03_reg[7]  ( .D(N89), .CP(clk), .Q(sa03[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][4]  ( .D(\u0/N244 ), .CP(clk), .Q(w3[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][10]  ( .D(\u0/N250 ), .CP(clk), .Q(w3[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][25]  ( .D(\u0/N265 ), .CP(clk), .Q(w3[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][7]  ( .D(\u0/N247 ), .CP(clk), .Q(w3[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][29]  ( .D(\u0/N269 ), .CP(clk), .Q(w3[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][31]  ( .D(\u0/N271 ), .CP(clk), .Q(w3[31]) );
  HS65_LL_DFPQX4 \sa20_reg[5]  ( .D(N247), .CP(clk), .Q(sa20[5]) );
  HS65_LL_DFPQX4 \sa11_reg[6]  ( .D(N200), .CP(clk), .Q(sa11[6]) );
  HS65_LL_DFPQX4 \sa21_reg[3]  ( .D(N181), .CP(clk), .Q(sa21[3]) );
  HS65_LL_DFPQX4 \sa20_reg[0]  ( .D(N242), .CP(clk), .Q(sa20[0]) );
  HS65_LL_DFPQX4 \sa30_reg[5]  ( .D(N231), .CP(clk), .Q(sa30[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][6]  ( .D(\u0/N246 ), .CP(clk), .Q(w3[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][26]  ( .D(\u0/N266 ), .CP(clk), .Q(w3[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][27]  ( .D(\u0/N267 ), .CP(clk), .Q(w3[27]) );
  HS65_LL_DFPQX4 \sa10_reg[5]  ( .D(N263), .CP(clk), .Q(sa10[5]) );
  HS65_LL_DFPQX4 \sa12_reg[6]  ( .D(N136), .CP(clk), .Q(sa12[6]) );
  HS65_LL_DFPQX4 \sa12_reg[1]  ( .D(N131), .CP(clk), .Q(sa12[1]) );
  HS65_LL_DFPQX4 \sa13_reg[6]  ( .D(N72), .CP(clk), .Q(sa13[6]) );
  HS65_LL_DFPQX4 \sa23_reg[7]  ( .D(N57), .CP(clk), .Q(sa23[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][28]  ( .D(\u0/N268 ), .CP(clk), .Q(w3[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][30]  ( .D(\u0/N270 ), .CP(clk), .Q(w3[30]) );
  HS65_LL_DFPQX4 \sa13_reg[7]  ( .D(N73), .CP(clk), .Q(sa13[7]) );
  HS65_LL_DFPQX4 \sa30_reg[3]  ( .D(N229), .CP(clk), .Q(sa30[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][24]  ( .D(\u0/N264 ), .CP(clk), .Q(w3[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][9]  ( .D(\u0/N249 ), .CP(clk), .Q(w3[9]) );
  HS65_LL_DFPQX4 \sa11_reg[1]  ( .D(N195), .CP(clk), .Q(sa11[1]) );
  HS65_LL_DFPQX4 \sa23_reg[5]  ( .D(N55), .CP(clk), .Q(sa23[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][3]  ( .D(\u0/N243 ), .CP(clk), .Q(w3[3]) );
  HS65_LL_DFPQX4 \sa00_reg[7]  ( .D(N281), .CP(clk), .Q(sa00[7]) );
  HS65_LL_DFPQX4 \sa10_reg[6]  ( .D(N264), .CP(clk), .Q(sa10[6]) );
  HS65_LL_DFPQX4 \sa21_reg[5]  ( .D(N183), .CP(clk), .Q(sa21[5]) );
  HS65_LL_DFPQX4 \sa12_reg[7]  ( .D(N137), .CP(clk), .Q(sa12[7]) );
  HS65_LL_DFPQX4 \sa32_reg[1]  ( .D(N99), .CP(clk), .Q(sa32[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][16]  ( .D(\u0/N256 ), .CP(clk), .Q(w3[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][0]  ( .D(\u0/N240 ), .CP(clk), .Q(w3[0]) );
  HS65_LL_DFPQX4 \sa02_reg[1]  ( .D(N147), .CP(clk), .Q(sa02[1]) );
  HS65_LL_DFPQX4 \sa12_reg[5]  ( .D(N135), .CP(clk), .Q(sa12[5]) );
  HS65_LL_DFPQX4 \sa02_reg[7]  ( .D(N153), .CP(clk), .Q(sa02[7]) );
  HS65_LL_DFPQX4 \sa02_reg[5]  ( .D(N151), .CP(clk), .Q(sa02[5]) );
  HS65_LL_DFPQX4 \sa23_reg[1]  ( .D(N51), .CP(clk), .Q(sa23[1]) );
  HS65_LL_DFPQX4 \sa11_reg[5]  ( .D(N199), .CP(clk), .Q(sa11[5]) );
  HS65_LL_DFPQX4 \sa10_reg[7]  ( .D(N265), .CP(clk), .Q(sa10[7]) );
  HS65_LL_DFPQX4 \sa01_reg[7]  ( .D(N217), .CP(clk), .Q(sa01[7]) );
  HS65_LL_DFPQX4 \sa33_reg[7]  ( .D(N41), .CP(clk), .Q(sa33[7]) );
  HS65_LL_DFPQX4 \sa20_reg[6]  ( .D(N248), .CP(clk), .Q(sa20[6]) );
  HS65_LL_DFPQX4 \sa21_reg[1]  ( .D(N179), .CP(clk), .Q(sa21[1]) );
  HS65_LL_DFPQX4 \sa00_reg[1]  ( .D(N275), .CP(clk), .Q(sa00[1]) );
  HS65_LL_DFPQX4 \sa21_reg[6]  ( .D(N184), .CP(clk), .Q(sa21[6]) );
  HS65_LL_DFPQX4 \sa31_reg[5]  ( .D(N167), .CP(clk), .Q(sa31[5]) );
  HS65_LL_DFPQX4 \sa03_reg[6]  ( .D(N88), .CP(clk), .Q(sa03[6]) );
  HS65_LL_DFPQX4 \sa03_reg[1]  ( .D(N83), .CP(clk), .Q(sa03[1]) );
  HS65_LL_DFPQX4 \sa31_reg[6]  ( .D(N168), .CP(clk), .Q(sa31[6]) );
  HS65_LL_DFPQX4 \sa31_reg[1]  ( .D(N163), .CP(clk), .Q(sa31[1]) );
  HS65_LL_OAI21X2 U13 ( .A(n3), .B(n7668), .C(n2), .Z(n7) );
  HS65_LL_AO312X4 U19 ( .A(n7665), .B(n8), .C(n7668), .D(dcnt[1]), .E(n7), .F(
        n6), .Z(n7670) );
  HS65_LL_OAI21X2 U21 ( .A(dcnt[0]), .B(n11), .C(n10), .Z(n7672) );
  HS65_LL_CB4I1X4 U20 ( .A(dcnt[3]), .B(n9), .C(n15842), .D(rst), .Z(n7671) );
  HS65_LL_NAND2X2 U6 ( .A(rst), .B(n15844), .Z(n3) );
  HS65_LL_IVX2 U11 ( .A(n8), .Z(n11) );
  HS65_LL_NAND3X2 U12 ( .A(rst), .B(n15843), .C(n11), .Z(n2) );
  HS65_LL_NAND2X2 U17 ( .A(n15842), .B(rst), .Z(n10) );
  HS65_LL_IVX2 U18 ( .A(n10), .Z(n6) );
  HS65_LL_NAND2X2 U8 ( .A(n1), .B(n8), .Z(n9) );
  HS65_LL_IVX2 U9 ( .A(n3), .Z(n4) );
  HS65_LL_CBI4I1X3 U14 ( .A(dcnt[1]), .B(n4), .C(n7), .D(dcnt[2]), .Z(n5) );
  HS65_LL_NAND2X2 U15 ( .A(n9), .B(n5), .Z(n7669) );
  HS65_LL_AOI12X2 U7 ( .A(n1), .B(n7664), .C(n3), .Z(n8) );
  HS65_LL_DFPHQX4 \text_in_r_reg[126]  ( .D(text_in[126]), .E(n7678), .CP(clk), 
        .Q(text_in_r[126]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[125]  ( .D(text_in[125]), .E(n15783), .CP(clk), .Q(text_in_r[125]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[124]  ( .D(text_in[124]), .E(n7678), .CP(clk), 
        .Q(text_in_r[124]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[123]  ( .D(text_in[123]), .E(n7677), .CP(clk), 
        .Q(text_in_r[123]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[122]  ( .D(text_in[122]), .E(n7676), .CP(clk), 
        .Q(text_in_r[122]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[121]  ( .D(text_in[121]), .E(n7675), .CP(clk), 
        .Q(text_in_r[121]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[120]  ( .D(text_in[120]), .E(n7674), .CP(clk), 
        .Q(text_in_r[120]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[119]  ( .D(text_in[119]), .E(n7673), .CP(clk), 
        .Q(text_in_r[119]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[118]  ( .D(text_in[118]), .E(n7675), .CP(clk), 
        .Q(text_in_r[118]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[117]  ( .D(text_in[117]), .E(n15783), .CP(clk), .Q(text_in_r[117]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[116]  ( .D(text_in[116]), .E(n7678), .CP(clk), 
        .Q(text_in_r[116]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[115]  ( .D(text_in[115]), .E(n7677), .CP(clk), 
        .Q(text_in_r[115]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[114]  ( .D(text_in[114]), .E(n7676), .CP(clk), 
        .Q(text_in_r[114]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[113]  ( .D(text_in[113]), .E(n7675), .CP(clk), 
        .Q(text_in_r[113]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[112]  ( .D(text_in[112]), .E(n7674), .CP(clk), 
        .Q(text_in_r[112]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[111]  ( .D(text_in[111]), .E(n7673), .CP(clk), 
        .Q(text_in_r[111]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[110]  ( .D(text_in[110]), .E(n7673), .CP(clk), 
        .Q(text_in_r[110]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[109]  ( .D(text_in[109]), .E(n15783), .CP(clk), .Q(text_in_r[109]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[108]  ( .D(text_in[108]), .E(n7678), .CP(clk), 
        .Q(text_in_r[108]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[107]  ( .D(text_in[107]), .E(n7677), .CP(clk), 
        .Q(text_in_r[107]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[106]  ( .D(text_in[106]), .E(n7676), .CP(clk), 
        .Q(text_in_r[106]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[105]  ( .D(text_in[105]), .E(n7675), .CP(clk), 
        .Q(text_in_r[105]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[104]  ( .D(text_in[104]), .E(n7674), .CP(clk), 
        .Q(text_in_r[104]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[103]  ( .D(text_in[103]), .E(n7673), .CP(clk), 
        .Q(text_in_r[103]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[102]  ( .D(text_in[102]), .E(n7674), .CP(clk), 
        .Q(text_in_r[102]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[101]  ( .D(text_in[101]), .E(n15839), .CP(clk), .Q(text_in_r[101]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[100]  ( .D(text_in[100]), .E(n7678), .CP(clk), 
        .Q(text_in_r[100]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[99]  ( .D(text_in[99]), .E(n7677), .CP(clk), 
        .Q(text_in_r[99]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[72]  ( .D(text_in[72]), .E(n7676), .CP(clk), 
        .Q(text_in_r[72]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[71]  ( .D(text_in[71]), .E(n7675), .CP(clk), 
        .Q(text_in_r[71]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[62]  ( .D(text_in[62]), .E(n7674), .CP(clk), 
        .Q(text_in_r[62]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[61]  ( .D(text_in[61]), .E(n7673), .CP(clk), 
        .Q(text_in_r[61]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[38]  ( .D(text_in[38]), .E(n7675), .CP(clk), 
        .Q(text_in_r[38]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[36]  ( .D(text_in[36]), .E(n15839), .CP(clk), 
        .Q(text_in_r[36]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[31]  ( .D(text_in[31]), .E(n7678), .CP(clk), 
        .Q(text_in_r[31]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[11]  ( .D(text_in[11]), .E(n7677), .CP(clk), 
        .Q(text_in_r[11]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[98]  ( .D(text_in[98]), .E(n7676), .CP(clk), 
        .Q(text_in_r[98]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[97]  ( .D(text_in[97]), .E(n7675), .CP(clk), 
        .Q(text_in_r[97]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[96]  ( .D(text_in[96]), .E(n7674), .CP(clk), 
        .Q(text_in_r[96]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[95]  ( .D(text_in[95]), .E(n7673), .CP(clk), 
        .Q(text_in_r[95]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[94]  ( .D(text_in[94]), .E(n7676), .CP(clk), 
        .Q(text_in_r[94]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[93]  ( .D(text_in[93]), .E(n15839), .CP(clk), 
        .Q(text_in_r[93]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[92]  ( .D(text_in[92]), .E(n7678), .CP(clk), 
        .Q(text_in_r[92]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[91]  ( .D(text_in[91]), .E(n7677), .CP(clk), 
        .Q(text_in_r[91]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[90]  ( .D(text_in[90]), .E(n7676), .CP(clk), 
        .Q(text_in_r[90]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[89]  ( .D(text_in[89]), .E(n7675), .CP(clk), 
        .Q(text_in_r[89]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[88]  ( .D(text_in[88]), .E(n7674), .CP(clk), 
        .Q(text_in_r[88]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[87]  ( .D(text_in[87]), .E(n7673), .CP(clk), 
        .Q(text_in_r[87]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[86]  ( .D(text_in[86]), .E(n7677), .CP(clk), 
        .Q(text_in_r[86]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[85]  ( .D(text_in[85]), .E(n15839), .CP(clk), 
        .Q(text_in_r[85]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[84]  ( .D(text_in[84]), .E(n7678), .CP(clk), 
        .Q(text_in_r[84]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[73]  ( .D(text_in[73]), .E(n7677), .CP(clk), 
        .Q(text_in_r[73]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[58]  ( .D(text_in[58]), .E(n7676), .CP(clk), 
        .Q(text_in_r[58]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[57]  ( .D(text_in[57]), .E(n7675), .CP(clk), 
        .Q(text_in_r[57]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[49]  ( .D(text_in[49]), .E(n7674), .CP(clk), 
        .Q(text_in_r[49]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[127]  ( .D(text_in[127]), .E(n7673), .CP(clk), 
        .Q(text_in_r[127]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[83]  ( .D(text_in[83]), .E(n7678), .CP(clk), 
        .Q(text_in_r[83]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[82]  ( .D(text_in[82]), .E(n15839), .CP(clk), 
        .Q(text_in_r[82]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[81]  ( .D(text_in[81]), .E(n7678), .CP(clk), 
        .Q(text_in_r[81]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[80]  ( .D(text_in[80]), .E(n7677), .CP(clk), 
        .Q(text_in_r[80]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[79]  ( .D(text_in[79]), .E(n7676), .CP(clk), 
        .Q(text_in_r[79]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[78]  ( .D(text_in[78]), .E(n7675), .CP(clk), 
        .Q(text_in_r[78]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[77]  ( .D(text_in[77]), .E(n7674), .CP(clk), 
        .Q(text_in_r[77]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[76]  ( .D(text_in[76]), .E(n7673), .CP(clk), 
        .Q(text_in_r[76]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[75]  ( .D(text_in[75]), .E(n7676), .CP(clk), 
        .Q(text_in_r[75]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[74]  ( .D(text_in[74]), .E(n7673), .CP(clk), 
        .Q(text_in_r[74]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[70]  ( .D(text_in[70]), .E(n7678), .CP(clk), 
        .Q(text_in_r[70]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[69]  ( .D(text_in[69]), .E(n7677), .CP(clk), 
        .Q(text_in_r[69]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[68]  ( .D(text_in[68]), .E(n7676), .CP(clk), 
        .Q(text_in_r[68]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[67]  ( .D(text_in[67]), .E(n7675), .CP(clk), 
        .Q(text_in_r[67]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[65]  ( .D(text_in[65]), .E(n7674), .CP(clk), 
        .Q(text_in_r[65]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[63]  ( .D(text_in[63]), .E(n7673), .CP(clk), 
        .Q(text_in_r[63]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[60]  ( .D(text_in[60]), .E(n7673), .CP(clk), 
        .Q(text_in_r[60]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[56]  ( .D(text_in[56]), .E(n7674), .CP(clk), 
        .Q(text_in_r[56]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[55]  ( .D(text_in[55]), .E(n7678), .CP(clk), 
        .Q(text_in_r[55]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[53]  ( .D(text_in[53]), .E(n7677), .CP(clk), 
        .Q(text_in_r[53]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[52]  ( .D(text_in[52]), .E(n7676), .CP(clk), 
        .Q(text_in_r[52]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[51]  ( .D(text_in[51]), .E(n7675), .CP(clk), 
        .Q(text_in_r[51]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[48]  ( .D(text_in[48]), .E(n7674), .CP(clk), 
        .Q(text_in_r[48]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[46]  ( .D(text_in[46]), .E(n7673), .CP(clk), 
        .Q(text_in_r[46]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[42]  ( .D(text_in[42]), .E(n7674), .CP(clk), 
        .Q(text_in_r[42]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[40]  ( .D(text_in[40]), .E(n7675), .CP(clk), 
        .Q(text_in_r[40]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[34]  ( .D(text_in[34]), .E(n7678), .CP(clk), 
        .Q(text_in_r[34]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[33]  ( .D(text_in[33]), .E(n7677), .CP(clk), 
        .Q(text_in_r[33]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[32]  ( .D(text_in[32]), .E(n7676), .CP(clk), 
        .Q(text_in_r[32]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[30]  ( .D(text_in[30]), .E(n7675), .CP(clk), 
        .Q(text_in_r[30]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[29]  ( .D(text_in[29]), .E(n7674), .CP(clk), 
        .Q(text_in_r[29]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[28]  ( .D(text_in[28]), .E(n7673), .CP(clk), 
        .Q(text_in_r[28]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[27]  ( .D(text_in[27]), .E(n7675), .CP(clk), 
        .Q(text_in_r[27]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[26]  ( .D(text_in[26]), .E(n7676), .CP(clk), 
        .Q(text_in_r[26]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[25]  ( .D(text_in[25]), .E(n7678), .CP(clk), 
        .Q(text_in_r[25]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[24]  ( .D(text_in[24]), .E(n7677), .CP(clk), 
        .Q(text_in_r[24]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[23]  ( .D(text_in[23]), .E(n7676), .CP(clk), 
        .Q(text_in_r[23]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[22]  ( .D(text_in[22]), .E(n7675), .CP(clk), 
        .Q(text_in_r[22]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[21]  ( .D(text_in[21]), .E(n7674), .CP(clk), 
        .Q(text_in_r[21]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[20]  ( .D(text_in[20]), .E(n7673), .CP(clk), 
        .Q(text_in_r[20]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[19]  ( .D(text_in[19]), .E(n7676), .CP(clk), 
        .Q(text_in_r[19]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[18]  ( .D(text_in[18]), .E(n7677), .CP(clk), 
        .Q(text_in_r[18]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[17]  ( .D(text_in[17]), .E(n7678), .CP(clk), 
        .Q(text_in_r[17]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[16]  ( .D(text_in[16]), .E(n7677), .CP(clk), 
        .Q(text_in_r[16]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[15]  ( .D(text_in[15]), .E(n7676), .CP(clk), 
        .Q(text_in_r[15]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[14]  ( .D(text_in[14]), .E(n7675), .CP(clk), 
        .Q(text_in_r[14]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[13]  ( .D(text_in[13]), .E(n7674), .CP(clk), 
        .Q(text_in_r[13]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[12]  ( .D(text_in[12]), .E(n7673), .CP(clk), 
        .Q(text_in_r[12]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[10]  ( .D(text_in[10]), .E(n7677), .CP(clk), 
        .Q(text_in_r[10]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[9]  ( .D(text_in[9]), .E(n7674), .CP(clk), 
        .Q(text_in_r[9]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[8]  ( .D(text_in[8]), .E(n7678), .CP(clk), 
        .Q(text_in_r[8]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[7]  ( .D(text_in[7]), .E(n7677), .CP(clk), 
        .Q(text_in_r[7]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[6]  ( .D(text_in[6]), .E(n7676), .CP(clk), 
        .Q(text_in_r[6]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[5]  ( .D(text_in[5]), .E(n7675), .CP(clk), 
        .Q(text_in_r[5]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[4]  ( .D(text_in[4]), .E(n7674), .CP(clk), 
        .Q(text_in_r[4]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[3]  ( .D(text_in[3]), .E(n7673), .CP(clk), 
        .Q(text_in_r[3]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[2]  ( .D(text_in[2]), .E(n7677), .CP(clk), 
        .Q(text_in_r[2]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[1]  ( .D(text_in[1]), .E(n7673), .CP(clk), 
        .Q(text_in_r[1]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[0]  ( .D(text_in[0]), .E(n7678), .CP(clk), 
        .Q(text_in_r[0]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[66]  ( .D(text_in[66]), .E(n7677), .CP(clk), 
        .Q(text_in_r[66]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[64]  ( .D(text_in[64]), .E(n7676), .CP(clk), 
        .Q(text_in_r[64]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[59]  ( .D(text_in[59]), .E(n7675), .CP(clk), 
        .Q(text_in_r[59]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[54]  ( .D(text_in[54]), .E(n7674), .CP(clk), 
        .Q(text_in_r[54]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[44]  ( .D(text_in[44]), .E(n7673), .CP(clk), 
        .Q(text_in_r[44]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[50]  ( .D(text_in[50]), .E(n7678), .CP(clk), 
        .Q(text_in_r[50]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[47]  ( .D(text_in[47]), .E(n7678), .CP(clk), 
        .Q(text_in_r[47]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[45]  ( .D(text_in[45]), .E(n7678), .CP(clk), 
        .Q(text_in_r[45]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[43]  ( .D(text_in[43]), .E(n7677), .CP(clk), 
        .Q(text_in_r[43]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[41]  ( .D(text_in[41]), .E(n7676), .CP(clk), 
        .Q(text_in_r[41]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[39]  ( .D(text_in[39]), .E(n7675), .CP(clk), 
        .Q(text_in_r[39]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[37]  ( .D(text_in[37]), .E(n7674), .CP(clk), 
        .Q(text_in_r[37]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[35]  ( .D(text_in[35]), .E(n7673), .CP(clk), 
        .Q(text_in_r[35]) );
  HS65_LLS_DFPQX18 \text_out_reg[105]  ( .D(N448), .CP(clk), .Q(text_out[105])
         );
  HS65_LLS_DFPQX18 \text_out_reg[61]  ( .D(N396), .CP(clk), .Q(text_out[61])
         );
  HS65_LLS_DFPQX18 \text_out_reg[1]  ( .D(N504), .CP(clk), .Q(text_out[1]) );
  HS65_LLS_DFPQX18 done_reg ( .D(N23), .CP(clk), .Q(done) );
  HS65_LLS_DFPQX18 \text_out_reg[65]  ( .D(N488), .CP(clk), .Q(text_out[65])
         );
  HS65_LLS_DFPQX18 \text_out_reg[81]  ( .D(N424), .CP(clk), .Q(text_out[81])
         );
  HS65_LLS_DFPQX18 \text_out_reg[33]  ( .D(N496), .CP(clk), .Q(text_out[33])
         );
  HS65_LLS_DFPQX18 \text_out_reg[111]  ( .D(N442), .CP(clk), .Q(text_out[111])
         );
  HS65_LLS_DFPQX18 \text_out_reg[110]  ( .D(N443), .CP(clk), .Q(text_out[110])
         );
  HS65_LLS_DFPQX18 \text_out_reg[9]  ( .D(N472), .CP(clk), .Q(text_out[9]) );
  HS65_LLS_DFPQX18 \text_out_reg[113]  ( .D(N416), .CP(clk), .Q(text_out[113])
         );
  HS65_LLS_DFPQX18 \text_out_reg[89]  ( .D(N392), .CP(clk), .Q(text_out[89])
         );
  HS65_LLS_DFPQX18 \text_out_reg[80]  ( .D(N425), .CP(clk), .Q(text_out[80])
         );
  HS65_LLS_DFPQX18 \text_out_reg[50]  ( .D(N431), .CP(clk), .Q(text_out[50])
         );
  HS65_LLS_DFPQX18 \text_out_reg[60]  ( .D(N397), .CP(clk), .Q(text_out[60])
         );
  HS65_LLS_DFPQX18 \text_out_reg[10]  ( .D(N471), .CP(clk), .Q(text_out[10])
         );
  HS65_LLS_DFPQX18 \text_out_reg[43]  ( .D(N462), .CP(clk), .Q(text_out[43])
         );
  HS65_LLS_DFPQX18 \text_out_reg[121]  ( .D(N384), .CP(clk), .Q(text_out[121])
         );
  HS65_LLS_DFPQX18 \text_out_reg[44]  ( .D(N461), .CP(clk), .Q(text_out[44])
         );
  HS65_LLS_DFPQX18 \text_out_reg[117]  ( .D(N412), .CP(clk), .Q(text_out[117])
         );
  HS65_LLS_DFPQX18 \text_out_reg[85]  ( .D(N420), .CP(clk), .Q(text_out[85])
         );
  HS65_LLS_DFPQX18 \text_out_reg[62]  ( .D(N395), .CP(clk), .Q(text_out[62])
         );
  HS65_LLS_DFPQX18 \text_out_reg[40]  ( .D(N465), .CP(clk), .Q(text_out[40])
         );
  HS65_LLS_DFPQX18 \text_out_reg[124]  ( .D(N381), .CP(clk), .Q(text_out[124])
         );
  HS65_LLS_DFPQX18 \text_out_reg[70]  ( .D(N483), .CP(clk), .Q(text_out[70])
         );
  HS65_LLS_DFPQX18 \text_out_reg[57]  ( .D(N400), .CP(clk), .Q(text_out[57])
         );
  HS65_LLS_DFPQX18 \text_out_reg[73]  ( .D(N456), .CP(clk), .Q(text_out[73])
         );
  HS65_LLS_DFPQX18 \text_out_reg[99]  ( .D(N478), .CP(clk), .Q(text_out[99])
         );
  HS65_LLS_DFPQX18 \text_out_reg[26]  ( .D(N407), .CP(clk), .Q(text_out[26])
         );
  HS65_LLS_DFPQX18 \text_out_reg[58]  ( .D(N399), .CP(clk), .Q(text_out[58])
         );
  HS65_LLS_DFPQX18 \text_out_reg[88]  ( .D(N393), .CP(clk), .Q(text_out[88])
         );
  HS65_LLS_DFPQX18 \text_out_reg[25]  ( .D(N408), .CP(clk), .Q(text_out[25])
         );
  HS65_LLS_DFPQX18 \text_out_reg[68]  ( .D(N485), .CP(clk), .Q(text_out[68])
         );
  HS65_LLS_DFPQX18 \text_out_reg[18]  ( .D(N439), .CP(clk), .Q(text_out[18])
         );
  HS65_LLS_DFPQX18 \text_out_reg[93]  ( .D(N388), .CP(clk), .Q(text_out[93])
         );
  HS65_LLS_DFPQX18 \text_out_reg[41]  ( .D(N464), .CP(clk), .Q(text_out[41])
         );
  HS65_LLS_DFPQX18 \text_out_reg[21]  ( .D(N436), .CP(clk), .Q(text_out[21])
         );
  HS65_LLS_DFPQX18 \text_out_reg[59]  ( .D(N398), .CP(clk), .Q(text_out[59])
         );
  HS65_LLS_DFPQX18 \text_out_reg[71]  ( .D(N482), .CP(clk), .Q(text_out[71])
         );
  HS65_LLS_DFPQX18 \text_out_reg[54]  ( .D(N427), .CP(clk), .Q(text_out[54])
         );
  HS65_LLS_DFPQX18 \text_out_reg[23]  ( .D(N434), .CP(clk), .Q(text_out[23])
         );
  HS65_LLS_DFPQX18 \text_out_reg[12]  ( .D(N469), .CP(clk), .Q(text_out[12])
         );
  HS65_LLS_DFPQX18 \text_out_reg[47]  ( .D(N458), .CP(clk), .Q(text_out[47])
         );
  HS65_LLS_DFPQX18 \text_out_reg[46]  ( .D(N459), .CP(clk), .Q(text_out[46])
         );
  HS65_LLS_DFPQX18 \text_out_reg[116]  ( .D(N413), .CP(clk), .Q(text_out[116])
         );
  HS65_LLS_DFPQX18 \text_out_reg[107]  ( .D(N446), .CP(clk), .Q(text_out[107])
         );
  HS65_LLS_DFPQX18 \text_out_reg[100]  ( .D(N477), .CP(clk), .Q(text_out[100])
         );
  HS65_LLS_DFPQX18 \text_out_reg[102]  ( .D(N475), .CP(clk), .Q(text_out[102])
         );
  HS65_LLS_DFPQX18 \text_out_reg[101]  ( .D(N476), .CP(clk), .Q(text_out[101])
         );
  HS65_LLS_DFPQX18 \text_out_reg[5]  ( .D(N500), .CP(clk), .Q(text_out[5]) );
  HS65_LLS_DFPQX18 \text_out_reg[3]  ( .D(N502), .CP(clk), .Q(text_out[3]) );
  HS65_LLS_DFPQX18 \text_out_reg[29]  ( .D(N404), .CP(clk), .Q(text_out[29])
         );
  HS65_LLS_DFPQX18 \text_out_reg[31]  ( .D(N402), .CP(clk), .Q(text_out[31])
         );
  HS65_LLS_DFPQX18 \text_out_reg[38]  ( .D(N491), .CP(clk), .Q(text_out[38])
         );
  HS65_LLS_DFPQX18 \text_out_reg[53]  ( .D(N428), .CP(clk), .Q(text_out[53])
         );
  HS65_LLS_DFPQX18 \text_out_reg[27]  ( .D(N406), .CP(clk), .Q(text_out[27])
         );
  HS65_LLS_DFPQX18 \text_out_reg[119]  ( .D(N410), .CP(clk), .Q(text_out[119])
         );
  HS65_LLS_DFPQX18 \text_out_reg[42]  ( .D(N463), .CP(clk), .Q(text_out[42])
         );
  HS65_LLS_DFPQX18 \text_out_reg[92]  ( .D(N389), .CP(clk), .Q(text_out[92])
         );
  HS65_LLS_DFPQX18 \text_out_reg[55]  ( .D(N426), .CP(clk), .Q(text_out[55])
         );
  HS65_LLS_DFPQX18 \text_out_reg[97]  ( .D(N480), .CP(clk), .Q(text_out[97])
         );
  HS65_LLS_DFPQX18 \text_out_reg[127]  ( .D(N378), .CP(clk), .Q(text_out[127])
         );
  HS65_LLS_DFPQX18 \text_out_reg[16]  ( .D(N441), .CP(clk), .Q(text_out[16])
         );
  HS65_LLS_DFPQX18 \text_out_reg[91]  ( .D(N390), .CP(clk), .Q(text_out[91])
         );
  HS65_LLS_DFPQX18 \text_out_reg[13]  ( .D(N468), .CP(clk), .Q(text_out[13])
         );
  HS65_LLS_DFPQX18 \text_out_reg[69]  ( .D(N484), .CP(clk), .Q(text_out[69])
         );
  HS65_LLS_DFPQX18 \text_out_reg[112]  ( .D(N417), .CP(clk), .Q(text_out[112])
         );
  HS65_LLS_DFPQX18 \text_out_reg[90]  ( .D(N391), .CP(clk), .Q(text_out[90])
         );
  HS65_LLS_DFPQX18 \text_out_reg[45]  ( .D(N460), .CP(clk), .Q(text_out[45])
         );
  HS65_LLS_DFPQX18 \text_out_reg[123]  ( .D(N382), .CP(clk), .Q(text_out[123])
         );
  HS65_LLS_DFPQX18 \text_out_reg[14]  ( .D(N467), .CP(clk), .Q(text_out[14])
         );
  HS65_LLS_DFPQX18 \text_out_reg[87]  ( .D(N418), .CP(clk), .Q(text_out[87])
         );
  HS65_LLS_DFPQX18 \text_out_reg[94]  ( .D(N387), .CP(clk), .Q(text_out[94])
         );
  HS65_LLS_DFPQX18 \text_out_reg[19]  ( .D(N438), .CP(clk), .Q(text_out[19])
         );
  HS65_LLS_DFPQX18 \text_out_reg[86]  ( .D(N419), .CP(clk), .Q(text_out[86])
         );
  HS65_LLS_DFPQX18 \text_out_reg[4]  ( .D(N501), .CP(clk), .Q(text_out[4]) );
  HS65_LLS_DFPQX18 \text_out_reg[115]  ( .D(N414), .CP(clk), .Q(text_out[115])
         );
  HS65_LLS_DFPQX18 \text_out_reg[51]  ( .D(N430), .CP(clk), .Q(text_out[51])
         );
  HS65_LLS_DFPQX18 \text_out_reg[36]  ( .D(N493), .CP(clk), .Q(text_out[36])
         );
  HS65_LLS_DFPQX18 \text_out_reg[82]  ( .D(N423), .CP(clk), .Q(text_out[82])
         );
  HS65_LLS_DFPQX18 \text_out_reg[34]  ( .D(N495), .CP(clk), .Q(text_out[34])
         );
  HS65_LLS_DFPQX18 \text_out_reg[77]  ( .D(N452), .CP(clk), .Q(text_out[77])
         );
  HS65_LLS_DFPQX18 \text_out_reg[15]  ( .D(N466), .CP(clk), .Q(text_out[15])
         );
  HS65_LLS_DFPQX18 \text_out_reg[52]  ( .D(N429), .CP(clk), .Q(text_out[52])
         );
  HS65_LLS_DFPQX18 \text_out_reg[72]  ( .D(N457), .CP(clk), .Q(text_out[72])
         );
  HS65_LLS_DFPQX18 \text_out_reg[103]  ( .D(N474), .CP(clk), .Q(text_out[103])
         );
  HS65_LLS_DFPQX18 \text_out_reg[48]  ( .D(N433), .CP(clk), .Q(text_out[48])
         );
  HS65_LLS_DFPQX18 \text_out_reg[106]  ( .D(N447), .CP(clk), .Q(text_out[106])
         );
  HS65_LLS_DFPQX18 \text_out_reg[83]  ( .D(N422), .CP(clk), .Q(text_out[83])
         );
  HS65_LLS_DFPQX18 \text_out_reg[108]  ( .D(N445), .CP(clk), .Q(text_out[108])
         );
  HS65_LLS_DFPQX18 \text_out_reg[96]  ( .D(N481), .CP(clk), .Q(text_out[96])
         );
  HS65_LLS_DFPQX18 \text_out_reg[84]  ( .D(N421), .CP(clk), .Q(text_out[84])
         );
  HS65_LLS_DFPQX18 \text_out_reg[49]  ( .D(N432), .CP(clk), .Q(text_out[49])
         );
  HS65_LLS_DFPQX18 \text_out_reg[75]  ( .D(N454), .CP(clk), .Q(text_out[75])
         );
  HS65_LLS_DFPQX18 \text_out_reg[17]  ( .D(N440), .CP(clk), .Q(text_out[17])
         );
  HS65_LLS_DFPQX18 \text_out_reg[79]  ( .D(N450), .CP(clk), .Q(text_out[79])
         );
  HS65_LLS_DFPQX18 \text_out_reg[7]  ( .D(N498), .CP(clk), .Q(text_out[7]) );
  HS65_LLS_DFPQX18 \text_out_reg[63]  ( .D(N394), .CP(clk), .Q(text_out[63])
         );
  HS65_LLS_DFPQX18 \text_out_reg[109]  ( .D(N444), .CP(clk), .Q(text_out[109])
         );
  HS65_LLS_DFPQX18 \text_out_reg[2]  ( .D(N503), .CP(clk), .Q(text_out[2]) );
  HS65_LLS_DFPQX18 \text_out_reg[104]  ( .D(N449), .CP(clk), .Q(text_out[104])
         );
  HS65_LLS_DFPQX18 \text_out_reg[66]  ( .D(N487), .CP(clk), .Q(text_out[66])
         );
  HS65_LLS_DFPQX18 \text_out_reg[22]  ( .D(N435), .CP(clk), .Q(text_out[22])
         );
  HS65_LLS_DFPQX18 \text_out_reg[126]  ( .D(N379), .CP(clk), .Q(text_out[126])
         );
  HS65_LLS_DFPQX18 \text_out_reg[125]  ( .D(N380), .CP(clk), .Q(text_out[125])
         );
  HS65_LLS_DFPQX18 \text_out_reg[98]  ( .D(N479), .CP(clk), .Q(text_out[98])
         );
  HS65_LLS_DFPQX18 \text_out_reg[95]  ( .D(N386), .CP(clk), .Q(text_out[95])
         );
  HS65_LLS_DFPQX18 \text_out_reg[0]  ( .D(N505), .CP(clk), .Q(text_out[0]) );
  HS65_LLS_DFPQX18 \text_out_reg[28]  ( .D(N405), .CP(clk), .Q(text_out[28])
         );
  HS65_LLS_DFPQX18 \text_out_reg[37]  ( .D(N492), .CP(clk), .Q(text_out[37])
         );
  HS65_LLS_DFPQX18 \text_out_reg[8]  ( .D(N473), .CP(clk), .Q(text_out[8]) );
  HS65_LLS_DFPQX18 \text_out_reg[120]  ( .D(N385), .CP(clk), .Q(text_out[120])
         );
  HS65_LLS_DFPQX18 \text_out_reg[6]  ( .D(N499), .CP(clk), .Q(text_out[6]) );
  HS65_LLS_DFPQX18 \text_out_reg[24]  ( .D(N409), .CP(clk), .Q(text_out[24])
         );
  HS65_LLS_DFPQX18 \text_out_reg[11]  ( .D(N470), .CP(clk), .Q(text_out[11])
         );
  HS65_LLS_DFPQX18 \text_out_reg[64]  ( .D(N489), .CP(clk), .Q(text_out[64])
         );
  HS65_LLS_DFPQX18 \text_out_reg[78]  ( .D(N451), .CP(clk), .Q(text_out[78])
         );
  HS65_LLS_DFPQX18 \text_out_reg[20]  ( .D(N437), .CP(clk), .Q(text_out[20])
         );
  HS65_LLS_DFPQX18 \text_out_reg[56]  ( .D(N401), .CP(clk), .Q(text_out[56])
         );
  HS65_LLS_DFPQX18 \text_out_reg[32]  ( .D(N497), .CP(clk), .Q(text_out[32])
         );
  HS65_LLS_DFPQX18 \text_out_reg[74]  ( .D(N455), .CP(clk), .Q(text_out[74])
         );
  HS65_LLS_DFPQX18 \text_out_reg[118]  ( .D(N411), .CP(clk), .Q(text_out[118])
         );
  HS65_LLS_DFPQX18 \text_out_reg[76]  ( .D(N453), .CP(clk), .Q(text_out[76])
         );
  HS65_LLS_DFPQX18 \text_out_reg[67]  ( .D(N486), .CP(clk), .Q(text_out[67])
         );
  HS65_LLS_DFPQX18 \text_out_reg[114]  ( .D(N415), .CP(clk), .Q(text_out[114])
         );
  HS65_LLS_DFPQX18 \text_out_reg[122]  ( .D(N383), .CP(clk), .Q(text_out[122])
         );
  HS65_LLS_DFPQX18 \text_out_reg[35]  ( .D(N494), .CP(clk), .Q(text_out[35])
         );
  HS65_LLS_DFPQX18 \text_out_reg[30]  ( .D(N403), .CP(clk), .Q(text_out[30])
         );
  HS65_LLS_DFPQX18 \text_out_reg[39]  ( .D(N490), .CP(clk), .Q(text_out[39])
         );
  HS65_LL_DFPQX4 ld_r_reg ( .D(n15842), .CP(clk), .Q(ld_r) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[24]  ( .D(\u0/r0/N70 ), .CP(clk), .Q(
        \u0/rcon [24]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[2]  ( .D(\u0/r0/N80 ), .CP(clk), .Q(
        \u0/r0/rcnt [2]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[30]  ( .D(\u0/r0/N76 ), .CP(clk), .Q(
        \u0/rcon [30]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[1]  ( .D(\u0/r0/N79 ), .CP(clk), .Q(
        \u0/r0/rcnt [1]) );
  HS65_LL_DFPQX4 \dcnt_reg[3]  ( .D(n7671), .CP(clk), .Q(dcnt[3]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[3]  ( .D(\u0/r0/N81 ), .CP(clk), .Q(
        \u0/r0/rcnt [3]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[0]  ( .D(\u0/r0/N78 ), .CP(clk), .Q(
        \u0/r0/rcnt [0]) );
  HS65_LL_DFPQX4 \dcnt_reg[0]  ( .D(n7672), .CP(clk), .Q(dcnt[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][21]  ( .D(\u0/N63 ), .CP(clk), .Q(w0[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][23]  ( .D(\u0/N65 ), .CP(clk), .Q(w0[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][18]  ( .D(\u0/N60 ), .CP(clk), .Q(w0[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][11]  ( .D(\u0/N53 ), .CP(clk), .Q(w0[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][20]  ( .D(\u0/N62 ), .CP(clk), .Q(w0[20]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[26]  ( .D(\u0/r0/N72 ), .CP(clk), .Q(
        \u0/rcon [26]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[31]  ( .D(\u0/r0/N77 ), .CP(clk), .Q(
        \u0/rcon [31]) );
  HS65_LL_DFPQX4 \dcnt_reg[1]  ( .D(n7670), .CP(clk), .Q(dcnt[1]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[29]  ( .D(\u0/r0/N75 ), .CP(clk), .Q(
        \u0/rcon [29]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][14]  ( .D(\u0/N56 ), .CP(clk), .Q(w0[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][17]  ( .D(\u0/N59 ), .CP(clk), .Q(w0[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][13]  ( .D(\u0/N55 ), .CP(clk), .Q(w0[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][5]  ( .D(\u0/N47 ), .CP(clk), .Q(w0[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][22]  ( .D(\u0/N64 ), .CP(clk), .Q(w0[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][8]  ( .D(\u0/N50 ), .CP(clk), .Q(w0[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][12]  ( .D(\u0/N54 ), .CP(clk), .Q(w0[12]) );
  HS65_LL_DFPQX4 \dcnt_reg[2]  ( .D(n7669), .CP(clk), .Q(dcnt[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][19]  ( .D(\u0/N61 ), .CP(clk), .Q(w0[19]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[27]  ( .D(\u0/r0/N73 ), .CP(clk), .Q(
        \u0/rcon [27]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][1]  ( .D(\u0/N43 ), .CP(clk), .Q(w0[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][15]  ( .D(\u0/N57 ), .CP(clk), .Q(w0[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][21]  ( .D(\u0/N129 ), .CP(clk), .Q(w1[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][18]  ( .D(\u0/N126 ), .CP(clk), .Q(w1[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][23]  ( .D(\u0/N131 ), .CP(clk), .Q(w1[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][11]  ( .D(\u0/N119 ), .CP(clk), .Q(w1[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][20]  ( .D(\u0/N128 ), .CP(clk), .Q(w1[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][2]  ( .D(\u0/N44 ), .CP(clk), .Q(w0[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][4]  ( .D(\u0/N46 ), .CP(clk), .Q(w0[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][7]  ( .D(\u0/N49 ), .CP(clk), .Q(w0[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][25]  ( .D(\u0/N67 ), .CP(clk), .Q(w0[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][31]  ( .D(\u0/N73 ), .CP(clk), .Q(w0[31]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[25]  ( .D(\u0/r0/N71 ), .CP(clk), .Q(
        \u0/rcon [25]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[28]  ( .D(\u0/r0/N74 ), .CP(clk), .Q(
        \u0/rcon [28]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][9]  ( .D(\u0/N51 ), .CP(clk), .Q(w0[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][0]  ( .D(\u0/N42 ), .CP(clk), .Q(w0[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][13]  ( .D(\u0/N121 ), .CP(clk), .Q(w1[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][18]  ( .D(\u0/N192 ), .CP(clk), .Q(w2[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][10]  ( .D(\u0/N52 ), .CP(clk), .Q(w0[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][14]  ( .D(\u0/N122 ), .CP(clk), .Q(w1[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][17]  ( .D(\u0/N125 ), .CP(clk), .Q(w1[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][12]  ( .D(\u0/N120 ), .CP(clk), .Q(w1[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][5]  ( .D(\u0/N113 ), .CP(clk), .Q(w1[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][19]  ( .D(\u0/N127 ), .CP(clk), .Q(w1[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][8]  ( .D(\u0/N116 ), .CP(clk), .Q(w1[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][22]  ( .D(\u0/N130 ), .CP(clk), .Q(w1[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][1]  ( .D(\u0/N109 ), .CP(clk), .Q(w1[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][3]  ( .D(\u0/N45 ), .CP(clk), .Q(w0[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][16]  ( .D(\u0/N58 ), .CP(clk), .Q(w0[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][15]  ( .D(\u0/N123 ), .CP(clk), .Q(w1[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][29]  ( .D(\u0/N71 ), .CP(clk), .Q(w0[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][28]  ( .D(\u0/N70 ), .CP(clk), .Q(w0[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][6]  ( .D(\u0/N48 ), .CP(clk), .Q(w0[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][21]  ( .D(\u0/N195 ), .CP(clk), .Q(w2[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][2]  ( .D(\u0/N110 ), .CP(clk), .Q(w1[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][25]  ( .D(\u0/N133 ), .CP(clk), .Q(w1[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][4]  ( .D(\u0/N112 ), .CP(clk), .Q(w1[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][7]  ( .D(\u0/N115 ), .CP(clk), .Q(w1[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][31]  ( .D(\u0/N139 ), .CP(clk), .Q(w1[31]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][13]  ( .D(\u0/N187 ), .CP(clk), .Q(w2[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][23]  ( .D(\u0/N197 ), .CP(clk), .Q(w2[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][21]  ( .D(\u0/N261 ), .CP(clk), .Q(w3[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][18]  ( .D(\u0/N258 ), .CP(clk), .Q(w3[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][9]  ( .D(\u0/N117 ), .CP(clk), .Q(w1[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][20]  ( .D(\u0/N194 ), .CP(clk), .Q(w2[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][11]  ( .D(\u0/N185 ), .CP(clk), .Q(w2[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][0]  ( .D(\u0/N108 ), .CP(clk), .Q(w1[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][27]  ( .D(\u0/N69 ), .CP(clk), .Q(w0[27]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][23]  ( .D(\u0/N263 ), .CP(clk), .Q(w3[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][10]  ( .D(\u0/N118 ), .CP(clk), .Q(w1[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][30]  ( .D(\u0/N72 ), .CP(clk), .Q(w0[30]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][20]  ( .D(\u0/N260 ), .CP(clk), .Q(w3[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][11]  ( .D(\u0/N251 ), .CP(clk), .Q(w3[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][29]  ( .D(\u0/N137 ), .CP(clk), .Q(w1[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][3]  ( .D(\u0/N111 ), .CP(clk), .Q(w1[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][16]  ( .D(\u0/N124 ), .CP(clk), .Q(w1[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][24]  ( .D(\u0/N66 ), .CP(clk), .Q(w0[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][5]  ( .D(\u0/N179 ), .CP(clk), .Q(w2[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][22]  ( .D(\u0/N196 ), .CP(clk), .Q(w2[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][8]  ( .D(\u0/N182 ), .CP(clk), .Q(w2[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][26]  ( .D(\u0/N68 ), .CP(clk), .Q(w0[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][14]  ( .D(\u0/N188 ), .CP(clk), .Q(w2[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][17]  ( .D(\u0/N191 ), .CP(clk), .Q(w2[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][25]  ( .D(\u0/N199 ), .CP(clk), .Q(w2[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][28]  ( .D(\u0/N136 ), .CP(clk), .Q(w1[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][12]  ( .D(\u0/N186 ), .CP(clk), .Q(w2[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][19]  ( .D(\u0/N193 ), .CP(clk), .Q(w2[19]) );
  HS65_LL_DFPQX4 \sa20_reg[7]  ( .D(N249), .CP(clk), .Q(sa20[7]) );
  HS65_LL_DFPQX4 \sa02_reg[6]  ( .D(N152), .CP(clk), .Q(sa02[6]) );
  HS65_LL_DFPQX4 \sa33_reg[2]  ( .D(N36), .CP(clk), .Q(sa33[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][1]  ( .D(\u0/N175 ), .CP(clk), .Q(w2[1]) );
  HS65_LL_DFPQX4 \sa01_reg[6]  ( .D(N216), .CP(clk), .Q(sa01[6]) );
  HS65_LL_DFPQX4 \sa01_reg[5]  ( .D(N215), .CP(clk), .Q(sa01[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][5]  ( .D(\u0/N245 ), .CP(clk), .Q(w3[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][22]  ( .D(\u0/N262 ), .CP(clk), .Q(w3[22]) );
  HS65_LL_DFPQX4 \sa02_reg[2]  ( .D(N148), .CP(clk), .Q(sa02[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][13]  ( .D(\u0/N253 ), .CP(clk), .Q(w3[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][8]  ( .D(\u0/N248 ), .CP(clk), .Q(w3[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][6]  ( .D(\u0/N114 ), .CP(clk), .Q(w1[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][15]  ( .D(\u0/N189 ), .CP(clk), .Q(w2[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][14]  ( .D(\u0/N254 ), .CP(clk), .Q(w3[14]) );
  HS65_LL_DFPQX4 \sa23_reg[2]  ( .D(N52), .CP(clk), .Q(sa23[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][17]  ( .D(\u0/N257 ), .CP(clk), .Q(w3[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][12]  ( .D(\u0/N252 ), .CP(clk), .Q(w3[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][19]  ( .D(\u0/N259 ), .CP(clk), .Q(w3[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][1]  ( .D(\u0/N241 ), .CP(clk), .Q(w3[1]) );
  HS65_LL_DFPQX4 \sa03_reg[5]  ( .D(N87), .CP(clk), .Q(sa03[5]) );
  HS65_LL_DFPQX4 \sa32_reg[2]  ( .D(N100), .CP(clk), .Q(sa32[2]) );
  HS65_LL_DFPQX4 \sa21_reg[2]  ( .D(N180), .CP(clk), .Q(sa21[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][2]  ( .D(\u0/N176 ), .CP(clk), .Q(w2[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][15]  ( .D(\u0/N255 ), .CP(clk), .Q(w3[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][7]  ( .D(\u0/N181 ), .CP(clk), .Q(w2[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][4]  ( .D(\u0/N178 ), .CP(clk), .Q(w2[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][29]  ( .D(\u0/N203 ), .CP(clk), .Q(w2[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][31]  ( .D(\u0/N205 ), .CP(clk), .Q(w2[31]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][27]  ( .D(\u0/N135 ), .CP(clk), .Q(w1[27]) );
  HS65_LL_DFPQX4 \sa21_reg[7]  ( .D(N185), .CP(clk), .Q(sa21[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][30]  ( .D(\u0/N138 ), .CP(clk), .Q(w1[30]) );
  HS65_LL_DFPQX4 \sa01_reg[1]  ( .D(N211), .CP(clk), .Q(sa01[1]) );
  HS65_LL_BFX4 U8072 ( .A(ld), .Z(n7673) );
  HS65_LL_BFX4 U8073 ( .A(ld), .Z(n7674) );
  HS65_LL_BFX4 U8074 ( .A(ld), .Z(n7675) );
  HS65_LL_BFX4 U8075 ( .A(ld), .Z(n7676) );
  HS65_LL_BFX4 U8076 ( .A(ld), .Z(n7677) );
  HS65_LL_BFX4 U8077 ( .A(ld), .Z(n7678) );
  HS65_LL_IVX4 U8078 ( .A(ld), .Z(n15108) );
  HS65_LL_BFX4 U8079 ( .A(n15108), .Z(n15844) );
  HS65_LL_BFX2 U8080 ( .A(n15844), .Z(n15806) );
  HS65_LL_IVX4 U8081 ( .A(n15806), .Z(n15842) );
  HS65_LL_NAND3X2 U8082 ( .A(\u0/r0/rcnt [2]), .B(\u0/r0/rcnt [0]), .C(
        \u0/r0/rcnt [1]), .Z(n14989) );
  HS65_LL_NAND2X2 U8083 ( .A(n15108), .B(n14989), .Z(\u0/r0/N70 ) );
  HS65_LL_NOR2X2 U8084 ( .A(dcnt[1]), .B(dcnt[2]), .Z(n15841) );
  HS65_LL_NOR4ABX2 U8085 ( .A(dcnt[0]), .B(n15841), .C(n15842), .D(dcnt[3]), 
        .Z(N23) );
  HS65_LL_NOR2X2 U8086 ( .A(\u0/r0/rcnt [3]), .B(n14989), .Z(n14999) );
  HS65_LL_AOI12X2 U8087 ( .A(\u0/r0/rcnt [3]), .B(n14989), .C(n14999), .Z(
        n14990) );
  HS65_LL_IVX2 U8088 ( .A(\u0/r0/rcnt [2]), .Z(n14992) );
  HS65_LL_NOR2X2 U8089 ( .A(n15842), .B(\u0/r0/rcnt [0]), .Z(\u0/r0/N78 ) );
  HS65_LL_IVX2 U8090 ( .A(\u0/r0/N78 ), .Z(n14991) );
  HS65_LL_NOR4ABX2 U8091 ( .A(\u0/r0/rcnt [1]), .B(n14990), .C(n14992), .D(
        n14991), .Z(\u0/r0/N77 ) );
  HS65_LL_IVX2 U8092 ( .A(w3[13]), .Z(n15707) );
  HS65_LL_IVX2 U8093 ( .A(w2[13]), .Z(n15618) );
  HS65_LL_IVX2 U8094 ( .A(w1[13]), .Z(n15362) );
  HS65_LL_IVX2 U8095 ( .A(w0[13]), .Z(n15541) );
  HS65_LL_IVX2 U8096 ( .A(w3[6]), .Z(n15737) );
  HS65_LL_NAND2X2 U8097 ( .A(w3[1]), .B(n15737), .Z(n9438) );
  HS65_LL_IVX2 U8098 ( .A(n9438), .Z(n9395) );
  HS65_LL_NAND2X2 U8099 ( .A(w3[7]), .B(n9395), .Z(n9262) );
  HS65_LL_IVX2 U8100 ( .A(w3[3]), .Z(n15517) );
  HS65_LL_NOR2X2 U8101 ( .A(n15517), .B(w3[0]), .Z(n7692) );
  HS65_LL_NAND2X2 U8102 ( .A(w3[5]), .B(n7692), .Z(n7705) );
  HS65_LL_NOR2X2 U8103 ( .A(n9262), .B(n7705), .Z(n9587) );
  HS65_LL_NOR2X2 U8104 ( .A(w3[7]), .B(n9438), .Z(n7714) );
  HS65_LL_IVX2 U8105 ( .A(n7714), .Z(n7701) );
  HS65_LL_NAND2X2 U8106 ( .A(n15517), .B(w3[0]), .Z(n7687) );
  HS65_LL_NOR2X2 U8107 ( .A(n7687), .B(w3[5]), .Z(n9244) );
  HS65_LL_IVX2 U8108 ( .A(n9244), .Z(n9436) );
  HS65_LL_NOR2X2 U8109 ( .A(n7701), .B(n9436), .Z(n9252) );
  HS65_LL_NOR2X2 U8110 ( .A(w3[1]), .B(n15737), .Z(n9793) );
  HS65_LL_NAND2X2 U8111 ( .A(w3[7]), .B(n9793), .Z(n7703) );
  HS65_LL_NOR2X2 U8112 ( .A(n7703), .B(n7705), .Z(n9276) );
  HS65_LL_NOR2X2 U8113 ( .A(n9252), .B(n9276), .Z(n9589) );
  HS65_LL_IVX2 U8114 ( .A(w3[5]), .Z(n15730) );
  HS65_LL_OR2X4 U8115 ( .A(n7687), .B(n15730), .Z(n7716) );
  HS65_LL_IVX2 U8116 ( .A(w3[7]), .Z(n15746) );
  HS65_LL_NAND3X2 U8117 ( .A(w3[6]), .B(w3[1]), .C(n15746), .Z(n7720) );
  HS65_LL_NOR2X2 U8118 ( .A(n7716), .B(n7720), .Z(n9250) );
  HS65_LL_IVX2 U8119 ( .A(n9250), .Z(n9387) );
  HS65_LL_NAND2X2 U8120 ( .A(n9589), .B(n9387), .Z(n9374) );
  HS65_LL_NAND2X2 U8121 ( .A(w3[6]), .B(w3[1]), .Z(n9392) );
  HS65_LL_NOR2X2 U8122 ( .A(n15746), .B(n9392), .Z(n9249) );
  HS65_LL_IVX2 U8123 ( .A(n7705), .Z(n9394) );
  HS65_LL_NAND2X2 U8124 ( .A(n9249), .B(n9394), .Z(n9273) );
  HS65_LL_NAND3X2 U8125 ( .A(w3[0]), .B(w3[3]), .C(w3[5]), .Z(n7690) );
  HS65_LL_NOR2X2 U8126 ( .A(n7690), .B(n7701), .Z(n9579) );
  HS65_LL_IVX2 U8127 ( .A(n7720), .Z(n7704) );
  HS65_LL_NAND2X2 U8128 ( .A(n7704), .B(n9394), .Z(n9625) );
  HS65_LL_IVX2 U8129 ( .A(n9625), .Z(n9440) );
  HS65_LL_NOR2X2 U8130 ( .A(n9579), .B(n9440), .Z(n9606) );
  HS65_LL_NAND2X2 U8131 ( .A(n15730), .B(n7692), .Z(n7707) );
  HS65_LL_NOR3X1 U8132 ( .A(w3[7]), .B(n9438), .C(n7707), .Z(n9576) );
  HS65_LL_IVX2 U8133 ( .A(n9576), .Z(n9413) );
  HS65_LL_NOR2X2 U8134 ( .A(n7716), .B(n7703), .Z(n9863) );
  HS65_LL_NOR2X2 U8135 ( .A(w3[6]), .B(w3[1]), .Z(n9245) );
  HS65_LL_NAND2X2 U8136 ( .A(n9245), .B(n15746), .Z(n7719) );
  HS65_LL_NOR2X2 U8137 ( .A(n7690), .B(n7719), .Z(n9638) );
  HS65_LL_NOR2X2 U8138 ( .A(n9863), .B(n9638), .Z(n9270) );
  HS65_LL_NOR3X1 U8139 ( .A(w3[0]), .B(w3[3]), .C(w3[5]), .Z(n7684) );
  HS65_LL_NAND2X2 U8140 ( .A(n9793), .B(n15746), .Z(n9437) );
  HS65_LL_IVX2 U8141 ( .A(n9437), .Z(n9380) );
  HS65_LL_NAND2X2 U8142 ( .A(n7684), .B(n9380), .Z(n9439) );
  HS65_LL_NAND2X2 U8143 ( .A(w3[7]), .B(n9245), .Z(n7706) );
  HS65_LL_NOR2X2 U8144 ( .A(n7687), .B(n7706), .Z(n9635) );
  HS65_LL_IVX2 U8145 ( .A(n9635), .Z(n9402) );
  HS65_LL_NOR2X2 U8146 ( .A(w3[5]), .B(n9402), .Z(n7680) );
  HS65_LL_NOR2X2 U8147 ( .A(w3[0]), .B(w3[3]), .Z(n7679) );
  HS65_LL_NAND2X2 U8148 ( .A(w3[5]), .B(n7679), .Z(n9391) );
  HS65_LL_NOR2X2 U8149 ( .A(n7720), .B(n9391), .Z(n9241) );
  HS65_LL_NOR3AX2 U8150 ( .A(n9439), .B(n7680), .C(n9241), .Z(n9853) );
  HS65_LL_IVX2 U8151 ( .A(n7706), .Z(n7717) );
  HS65_LL_NAND2X2 U8152 ( .A(n7684), .B(n7717), .Z(n9396) );
  HS65_LL_IVX2 U8153 ( .A(n9396), .Z(n9569) );
  HS65_LL_NOR2X2 U8154 ( .A(n9438), .B(n7716), .Z(n9238) );
  HS65_LL_NAND2X2 U8155 ( .A(w3[7]), .B(n9238), .Z(n9860) );
  HS65_LL_NAND2X2 U8156 ( .A(n7684), .B(n7704), .Z(n9798) );
  HS65_LL_NAND2X2 U8157 ( .A(n9860), .B(n9798), .Z(n9836) );
  HS65_LL_NOR3AX2 U8158 ( .A(n9853), .B(n9569), .C(n9836), .Z(n9259) );
  HS65_LL_IVX2 U8159 ( .A(n7684), .Z(n9261) );
  HS65_LL_NOR2X2 U8160 ( .A(n9261), .B(n7719), .Z(n9584) );
  HS65_LL_CBI4I6X2 U8161 ( .A(n7714), .B(n9245), .C(n9394), .D(n9584), .Z(
        n7681) );
  HS65_LL_NAND3X2 U8162 ( .A(n9270), .B(n9259), .C(n7681), .Z(n9458) );
  HS65_LL_NAND3X2 U8163 ( .A(w3[3]), .B(w3[0]), .C(n15730), .Z(n7702) );
  HS65_LL_NOR2X2 U8164 ( .A(n7719), .B(n7702), .Z(n9791) );
  HS65_LL_NAND2X2 U8165 ( .A(n7684), .B(n9249), .Z(n9582) );
  HS65_LL_IVX2 U8166 ( .A(n9582), .Z(n7713) );
  HS65_LL_NOR2X2 U8167 ( .A(n9791), .B(n7713), .Z(n9449) );
  HS65_LL_NOR2X2 U8168 ( .A(n7703), .B(n9391), .Z(n7715) );
  HS65_LL_NOR2X2 U8169 ( .A(n7690), .B(n9437), .Z(n9639) );
  HS65_LL_NAND2X2 U8170 ( .A(n9244), .B(n9380), .Z(n9378) );
  HS65_LL_NOR2AX3 U8171 ( .A(n9249), .B(n7716), .Z(n9450) );
  HS65_LL_IVX2 U8172 ( .A(n9450), .Z(n9409) );
  HS65_LL_NAND2X2 U8173 ( .A(n9378), .B(n9409), .Z(n9583) );
  HS65_LL_NOR3X1 U8174 ( .A(n7715), .B(n9639), .C(n9583), .Z(n9247) );
  HS65_LL_IVX2 U8175 ( .A(w3[0]), .Z(n15717) );
  HS65_LL_NOR3X1 U8176 ( .A(n15717), .B(n15517), .C(n7706), .Z(n9581) );
  HS65_LL_NAND2X2 U8177 ( .A(w3[5]), .B(n9581), .Z(n9411) );
  HS65_LL_NAND3X2 U8178 ( .A(n9449), .B(n9247), .C(n9411), .Z(n7682) );
  HS65_LL_NOR4ABX2 U8179 ( .A(n9606), .B(n9413), .C(n9458), .D(n7682), .Z(
        n7683) );
  HS65_LL_NAND4ABX3 U8180 ( .A(n9587), .B(n9374), .C(n9273), .D(n7683), .Z(
        n7729) );
  HS65_LL_NAND2X2 U8181 ( .A(w3[2]), .B(w3[4]), .Z(n9875) );
  HS65_LL_IVX2 U8182 ( .A(n9875), .Z(n9599) );
  HS65_LL_NOR2X2 U8183 ( .A(n7690), .B(n7720), .Z(n9375) );
  HS65_LL_NOR2X2 U8184 ( .A(n9639), .B(n9584), .Z(n7718) );
  HS65_LL_OR2X4 U8185 ( .A(n7703), .B(n9436), .Z(n9817) );
  HS65_LL_NAND3AX3 U8186 ( .A(n9375), .B(n7718), .C(n9817), .Z(n9573) );
  HS65_LL_IVX2 U8187 ( .A(n7702), .Z(n7698) );
  HS65_LL_NAND2X2 U8188 ( .A(n9245), .B(n7698), .Z(n9852) );
  HS65_LL_NOR2X2 U8189 ( .A(n15746), .B(n9852), .Z(n7699) );
  HS65_LL_NOR2X2 U8190 ( .A(n7716), .B(n9437), .Z(n9258) );
  HS65_LL_NOR2X2 U8191 ( .A(n9391), .B(n7706), .Z(n9605) );
  HS65_LL_NOR2X2 U8192 ( .A(n9258), .B(n9605), .Z(n9641) );
  HS65_LL_IVX2 U8193 ( .A(n9641), .Z(n9272) );
  HS65_LL_NOR2X2 U8194 ( .A(n9863), .B(n9272), .Z(n7711) );
  HS65_LL_NAND2X2 U8195 ( .A(n7714), .B(n7692), .Z(n9843) );
  HS65_LL_NOR2X2 U8196 ( .A(n9262), .B(n9436), .Z(n9603) );
  HS65_LL_NOR2X2 U8197 ( .A(n9250), .B(n9603), .Z(n9811) );
  HS65_LL_NOR2X2 U8198 ( .A(n7690), .B(n9262), .Z(n9455) );
  HS65_LL_NOR2X2 U8199 ( .A(n9262), .B(n7707), .Z(n9619) );
  HS65_LL_NOR3X1 U8200 ( .A(n9455), .B(n7715), .C(n9619), .Z(n7685) );
  HS65_LL_NAND2X2 U8201 ( .A(n7684), .B(n7714), .Z(n9799) );
  HS65_LL_NAND3X2 U8202 ( .A(n9811), .B(n7685), .C(n9799), .Z(n9264) );
  HS65_LL_NOR4ABX2 U8203 ( .A(n7711), .B(n9843), .C(n9579), .D(n9264), .Z(
        n7686) );
  HS65_LL_OAI21X2 U8204 ( .A(n7687), .B(n7719), .C(n7686), .Z(n9572) );
  HS65_LL_NOR2X2 U8205 ( .A(n7699), .B(n9572), .Z(n9408) );
  HS65_LL_NAND2X2 U8206 ( .A(w3[5]), .B(n9635), .Z(n9839) );
  HS65_LL_NOR2X2 U8207 ( .A(n9261), .B(n7703), .Z(n9239) );
  HS65_LL_IVX2 U8208 ( .A(n9587), .Z(n9404) );
  HS65_LL_NAND2X2 U8209 ( .A(n9244), .B(n9249), .Z(n9257) );
  HS65_LL_NAND2X2 U8210 ( .A(n9404), .B(n9257), .Z(n7688) );
  HS65_LL_NOR4ABX2 U8211 ( .A(n9798), .B(n9839), .C(n9239), .D(n7688), .Z(
        n7689) );
  HS65_LL_NAND4ABX3 U8212 ( .A(n9252), .B(n9638), .C(n9408), .D(n7689), .Z(
        n7697) );
  HS65_LL_IVX2 U8213 ( .A(n7690), .Z(n9792) );
  HS65_LL_NAND2X2 U8214 ( .A(n9792), .B(n9249), .Z(n9452) );
  HS65_LL_IVX2 U8215 ( .A(n9793), .Z(n7691) );
  HS65_LL_NOR2X2 U8216 ( .A(n7691), .B(n7707), .Z(n9627) );
  HS65_LL_NAND2X2 U8217 ( .A(w3[7]), .B(n9627), .Z(n9383) );
  HS65_LL_NAND2X2 U8218 ( .A(n9452), .B(n9383), .Z(n9568) );
  HS65_LL_NOR2X2 U8219 ( .A(w3[7]), .B(n7702), .Z(n7700) );
  HS65_LL_NAND2X2 U8220 ( .A(n9793), .B(n7700), .Z(n7722) );
  HS65_LL_IVX2 U8221 ( .A(n7722), .Z(n9240) );
  HS65_LL_NOR2X2 U8222 ( .A(n9262), .B(n9391), .Z(n9810) );
  HS65_LL_NOR2X2 U8223 ( .A(n9240), .B(n9810), .Z(n9255) );
  HS65_LL_IVX2 U8224 ( .A(n7707), .Z(n7723) );
  HS65_LL_NAND2X2 U8225 ( .A(n7723), .B(n9249), .Z(n9268) );
  HS65_LL_NAND2X2 U8226 ( .A(n9255), .B(n9268), .Z(n9795) );
  HS65_LL_IVX2 U8227 ( .A(n7719), .Z(n7693) );
  HS65_LL_NAND2X2 U8228 ( .A(n15746), .B(n9238), .Z(n9643) );
  HS65_LL_IVX2 U8229 ( .A(n9643), .Z(n9801) );
  HS65_LL_AOI12X2 U8230 ( .A(n7693), .B(n7692), .C(n9801), .Z(n9382) );
  HS65_LL_NAND2X2 U8231 ( .A(w3[1]), .B(n7700), .Z(n9263) );
  HS65_LL_NAND3X2 U8232 ( .A(n9382), .B(n9582), .C(n9263), .Z(n7694) );
  HS65_LL_NOR3X1 U8233 ( .A(n9568), .B(n9795), .C(n7694), .Z(n9868) );
  HS65_LL_IVX2 U8234 ( .A(n9262), .Z(n7695) );
  HS65_LL_NAND2X2 U8235 ( .A(n7695), .B(n7698), .Z(n9251) );
  HS65_LL_IVX2 U8236 ( .A(n9251), .Z(n7696) );
  HS65_LL_NOR2X2 U8237 ( .A(n9391), .B(n7719), .Z(n9618) );
  HS65_LL_NOR3X1 U8238 ( .A(n7696), .B(n9241), .C(n9618), .Z(n9632) );
  HS65_LL_NAND4ABX3 U8239 ( .A(n9573), .B(n7697), .C(n9868), .D(n9632), .Z(
        n7728) );
  HS65_LL_NOR2X2 U8240 ( .A(w3[2]), .B(w3[4]), .Z(n9873) );
  HS65_LL_NOR2X2 U8241 ( .A(n7701), .B(n7702), .Z(n9634) );
  HS65_LL_NOR3X1 U8242 ( .A(n9455), .B(n9634), .C(n9810), .Z(n9647) );
  HS65_LL_NAND2X2 U8243 ( .A(n9249), .B(n7698), .Z(n9405) );
  HS65_LL_IVX2 U8244 ( .A(n9405), .Z(n9377) );
  HS65_LL_IVX2 U8245 ( .A(n9257), .Z(n9809) );
  HS65_LL_NOR3X1 U8246 ( .A(n9377), .B(n9587), .C(n9809), .Z(n9797) );
  HS65_LL_AOI12X2 U8247 ( .A(n7723), .B(n9395), .C(n9375), .Z(n9280) );
  HS65_LL_NAND3X2 U8248 ( .A(n9797), .B(n9280), .C(n9396), .Z(n9626) );
  HS65_LL_NOR2X2 U8249 ( .A(n7699), .B(n9626), .Z(n9806) );
  HS65_LL_NAND3X2 U8250 ( .A(w3[6]), .B(w3[1]), .C(n7700), .Z(n9410) );
  HS65_LL_NOR3X1 U8251 ( .A(w3[0]), .B(w3[3]), .C(n7701), .Z(n9620) );
  HS65_LL_NAND2X2 U8252 ( .A(w3[5]), .B(n9620), .Z(n9414) );
  HS65_LL_IVX2 U8253 ( .A(n9414), .Z(n9454) );
  HS65_LL_NOR3AX2 U8254 ( .A(n9410), .B(n9579), .C(n9454), .Z(n9832) );
  HS65_LL_IVX2 U8255 ( .A(n9832), .Z(n9819) );
  HS65_LL_NOR2X2 U8256 ( .A(n7703), .B(n7702), .Z(n9447) );
  HS65_LL_NOR3X1 U8257 ( .A(n9447), .B(n9639), .C(n9239), .Z(n9435) );
  HS65_LL_IVX2 U8258 ( .A(n9435), .Z(n9393) );
  HS65_LL_NOR3X1 U8259 ( .A(n7713), .B(n9819), .C(n9393), .Z(n7709) );
  HS65_LL_NOR2X2 U8260 ( .A(n9437), .B(n7705), .Z(n9591) );
  HS65_LL_NAND2X2 U8261 ( .A(n7704), .B(n9244), .Z(n9425) );
  HS65_LL_NAND3X2 U8262 ( .A(n9817), .B(n9425), .C(n9273), .Z(n7712) );
  HS65_LL_NAND2X2 U8263 ( .A(n7704), .B(n7723), .Z(n9616) );
  HS65_LL_IVX2 U8264 ( .A(n9252), .Z(n9567) );
  HS65_LL_NOR2X2 U8265 ( .A(n7706), .B(n7705), .Z(n9577) );
  HS65_LL_NOR2X2 U8266 ( .A(n7707), .B(n7719), .Z(n9456) );
  HS65_LL_NOR4ABX2 U8267 ( .A(n9616), .B(n9567), .C(n9577), .D(n9456), .Z(
        n7708) );
  HS65_LL_NAND4ABX3 U8268 ( .A(n9591), .B(n7712), .C(n7708), .D(n9860), .Z(
        n9812) );
  HS65_LL_NOR4ABX2 U8269 ( .A(n9806), .B(n7709), .C(n9627), .D(n9812), .Z(
        n7710) );
  HS65_LL_NAND3X2 U8270 ( .A(n7711), .B(n9647), .C(n7710), .Z(n7727) );
  HS65_LL_IVX2 U8271 ( .A(w3[2]), .Z(n15723) );
  HS65_LL_NAND2X2 U8272 ( .A(w3[4]), .B(n15723), .Z(n9866) );
  HS65_LL_IVX2 U8273 ( .A(n9866), .Z(n9609) );
  HS65_LL_NAND3X2 U8274 ( .A(n9245), .B(n9394), .C(n15746), .Z(n9849) );
  HS65_LL_NAND2X2 U8275 ( .A(n9799), .B(n9849), .Z(n9434) );
  HS65_LL_NOR2X2 U8276 ( .A(n9434), .B(n7712), .Z(n9840) );
  HS65_LL_AOI12X2 U8277 ( .A(n9394), .B(n7714), .C(n7713), .Z(n9803) );
  HS65_LL_IVX2 U8278 ( .A(n7715), .Z(n9269) );
  HS65_LL_NAND2X2 U8279 ( .A(n9269), .B(n9251), .Z(n9833) );
  HS65_LL_NOR2X2 U8280 ( .A(n7716), .B(n7719), .Z(n9446) );
  HS65_LL_IVX2 U8281 ( .A(n9446), .Z(n9275) );
  HS65_LL_NAND2X2 U8282 ( .A(n7723), .B(n7717), .Z(n9574) );
  HS65_LL_NAND2X2 U8283 ( .A(n9275), .B(n9574), .Z(n9389) );
  HS65_LL_NOR4ABX2 U8284 ( .A(n7718), .B(n9803), .C(n9833), .D(n9389), .Z(
        n9631) );
  HS65_LL_NOR2X2 U8285 ( .A(n9436), .B(n7719), .Z(n9593) );
  HS65_LL_NOR2X2 U8286 ( .A(n9593), .B(n9456), .Z(n9277) );
  HS65_LL_AOI12X2 U8287 ( .A(n7720), .B(n7719), .C(n9391), .Z(n7721) );
  HS65_LL_NOR4ABX2 U8288 ( .A(n9631), .B(n9277), .C(n9576), .D(n7721), .Z(
        n9427) );
  HS65_LL_AND2X4 U8289 ( .A(n9616), .B(n9378), .Z(n9403) );
  HS65_LL_NAND2X2 U8290 ( .A(n7722), .B(n9414), .Z(n9850) );
  HS65_LL_NOR4ABX2 U8291 ( .A(n9403), .B(n9404), .C(n9447), .D(n9850), .Z(
        n7724) );
  HS65_LL_NAND2X2 U8292 ( .A(n7723), .B(n9380), .Z(n9430) );
  HS65_LL_IVX2 U8293 ( .A(n9430), .Z(n9578) );
  HS65_LL_NOR4ABX2 U8294 ( .A(n9647), .B(n7724), .C(n9578), .D(n9375), .Z(
        n7725) );
  HS65_LL_NAND3X2 U8295 ( .A(n9840), .B(n9427), .C(n7725), .Z(n7726) );
  HS65_LL_IVX2 U8296 ( .A(w3[4]), .Z(n15515) );
  HS65_LL_NAND2X2 U8297 ( .A(w3[2]), .B(n15515), .Z(n9854) );
  HS65_LL_IVX2 U8298 ( .A(n9854), .Z(n9461) );
  HS65_LL_MX41X4 U8299 ( .D0(n7729), .S0(n9599), .D1(n7728), .S1(n9873), .D2(
        n7727), .S2(n9609), .D3(n7726), .S3(n9461), .Z(n7730) );
  HS65_LL_MUXI21X2 U8300 ( .D0(w0[13]), .D1(n15541), .S0(n7730), .Z(n9749) );
  HS65_LL_MUXI21X2 U8301 ( .D0(n15362), .D1(w1[13]), .S0(n9749), .Z(n10086) );
  HS65_LL_MUXI21X2 U8302 ( .D0(n15618), .D1(w2[13]), .S0(n10086), .Z(n10404)
         );
  HS65_LL_IVX4 U8303 ( .A(n15806), .Z(n15783) );
  HS65_LL_MUX31X4 U8304 ( .D0(n15707), .D1(w3[13]), .D2(key[13]), .S0(n10404), 
        .S1(n15783), .Z(\u0/N253 ) );
  HS65_LL_IVX2 U8305 ( .A(w3[25]), .Z(n15250) );
  HS65_LL_IVX2 U8306 ( .A(w2[25]), .Z(n15193) );
  HS65_LL_IVX2 U8307 ( .A(w1[25]), .Z(n15136) );
  HS65_LL_IVX2 U8308 ( .A(w3[19]), .Z(n15341) );
  HS65_LL_NOR2X2 U8309 ( .A(w3[16]), .B(n15341), .Z(n8012) );
  HS65_LL_IVX2 U8310 ( .A(w3[21]), .Z(n15681) );
  HS65_LL_NAND2X2 U8311 ( .A(n8012), .B(n15681), .Z(n7761) );
  HS65_LL_IVX2 U8312 ( .A(w3[23]), .Z(n15691) );
  HS65_LL_IVX2 U8313 ( .A(w3[22]), .Z(n15687) );
  HS65_LL_NAND2X2 U8314 ( .A(w3[17]), .B(n15687), .Z(n15047) );
  HS65_LL_NOR2X2 U8315 ( .A(n15691), .B(n15047), .Z(n7754) );
  HS65_LL_IVX2 U8316 ( .A(n7754), .Z(n7762) );
  HS65_LL_NOR2X2 U8317 ( .A(n7761), .B(n7762), .Z(n10456) );
  HS65_LL_NAND2X2 U8318 ( .A(w3[17]), .B(w3[22]), .Z(n7733) );
  HS65_LL_NOR2X2 U8319 ( .A(w3[23]), .B(n7733), .Z(n7737) );
  HS65_LL_IVX2 U8320 ( .A(n7737), .Z(n7748) );
  HS65_LL_NOR2X2 U8321 ( .A(n7761), .B(n7748), .Z(n10484) );
  HS65_LL_NOR3X1 U8322 ( .A(w3[16]), .B(w3[19]), .C(n15681), .Z(n7752) );
  HS65_LL_IVX2 U8323 ( .A(n7752), .Z(n7746) );
  HS65_LL_NOR2X2 U8324 ( .A(n7762), .B(n7746), .Z(n10340) );
  HS65_LL_IVX2 U8325 ( .A(n10340), .Z(n10489) );
  HS65_LL_NOR3X1 U8326 ( .A(w3[17]), .B(w3[22]), .C(w3[23]), .Z(n8026) );
  HS65_LL_NAND2X2 U8327 ( .A(n8026), .B(n7752), .Z(n10446) );
  HS65_LL_NAND4ABX3 U8328 ( .A(n10456), .B(n10484), .C(n10489), .D(n10446), 
        .Z(n7772) );
  HS65_LL_IVX2 U8329 ( .A(w3[17]), .Z(n15344) );
  HS65_LL_NAND2X2 U8330 ( .A(w3[22]), .B(n15344), .Z(n10523) );
  HS65_LL_NAND3X2 U8331 ( .A(w3[16]), .B(w3[19]), .C(w3[21]), .Z(n10524) );
  HS65_LL_NOR3X1 U8332 ( .A(n15691), .B(n10523), .C(n10524), .Z(n10332) );
  HS65_LL_NOR2X2 U8333 ( .A(w3[23]), .B(n15047), .Z(n8023) );
  HS65_LL_IVX2 U8334 ( .A(n8023), .Z(n7740) );
  HS65_LL_NOR3X1 U8335 ( .A(w3[16]), .B(w3[19]), .C(n7740), .Z(n10352) );
  HS65_LL_IVX2 U8336 ( .A(w3[16]), .Z(n15671) );
  HS65_LL_NOR2X2 U8337 ( .A(w3[19]), .B(n15671), .Z(n7763) );
  HS65_LL_NAND2X2 U8338 ( .A(w3[21]), .B(n7763), .Z(n8018) );
  HS65_LL_NOR2X2 U8339 ( .A(w3[23]), .B(n10523), .Z(n7735) );
  HS65_LL_IVX2 U8340 ( .A(n7735), .Z(n8043) );
  HS65_LL_NOR2X2 U8341 ( .A(n8018), .B(n8043), .Z(n10496) );
  HS65_LL_NAND3X2 U8342 ( .A(w3[17]), .B(w3[22]), .C(w3[23]), .Z(n15048) );
  HS65_LL_NAND2X2 U8343 ( .A(w3[21]), .B(n8012), .Z(n15046) );
  HS65_LL_NOR2X2 U8344 ( .A(n15048), .B(n15046), .Z(n10443) );
  HS65_LL_NOR2X2 U8345 ( .A(n10496), .B(n10443), .Z(n10448) );
  HS65_LL_NAND2X2 U8346 ( .A(n7763), .B(n15681), .Z(n10322) );
  HS65_LL_NOR2X2 U8347 ( .A(n10322), .B(n8043), .Z(n10485) );
  HS65_LL_NAND2X2 U8348 ( .A(w3[16]), .B(w3[19]), .Z(n7734) );
  HS65_LL_NOR2X2 U8349 ( .A(w3[21]), .B(n7734), .Z(n10422) );
  HS65_LL_IVX2 U8350 ( .A(n10422), .Z(n8035) );
  HS65_LL_NOR2X2 U8351 ( .A(n15048), .B(n8035), .Z(n10459) );
  HS65_LL_NAND3X2 U8352 ( .A(w3[16]), .B(w3[21]), .C(n7737), .Z(n10344) );
  HS65_LL_NOR2X2 U8353 ( .A(n15691), .B(n10523), .Z(n7753) );
  HS65_LL_IVX2 U8354 ( .A(n7753), .Z(n8036) );
  HS65_LL_NOR2X2 U8355 ( .A(n8036), .B(n15046), .Z(n15056) );
  HS65_LL_NOR3X1 U8356 ( .A(w3[23]), .B(n15047), .C(n10322), .Z(n10376) );
  HS65_LL_NOR2X2 U8357 ( .A(n15056), .B(n10376), .Z(n10363) );
  HS65_LL_NAND2X2 U8358 ( .A(n10344), .B(n10363), .Z(n15067) );
  HS65_LL_NOR3X1 U8359 ( .A(n10485), .B(n10459), .C(n15067), .Z(n7731) );
  HS65_LL_NOR3X1 U8360 ( .A(w3[16]), .B(w3[19]), .C(w3[21]), .Z(n7751) );
  HS65_LL_NAND2X2 U8361 ( .A(n7751), .B(n7754), .Z(n10362) );
  HS65_LL_NAND3X2 U8362 ( .A(n10448), .B(n7731), .C(n10362), .Z(n10409) );
  HS65_LL_NOR3X1 U8363 ( .A(n10332), .B(n10352), .C(n10409), .Z(n10414) );
  HS65_LL_IVX2 U8364 ( .A(n15047), .Z(n10324) );
  HS65_LL_IVX2 U8365 ( .A(n8018), .Z(n7732) );
  HS65_LL_NAND2X2 U8366 ( .A(n10324), .B(n7732), .Z(n8020) );
  HS65_LL_NOR2X2 U8367 ( .A(n10524), .B(n7762), .Z(n10316) );
  HS65_LL_NOR3X1 U8368 ( .A(w3[23]), .B(n10523), .C(n7761), .Z(n10464) );
  HS65_LL_NOR3AX2 U8369 ( .A(n8020), .B(n10316), .C(n10464), .Z(n10442) );
  HS65_LL_NOR3X1 U8370 ( .A(w3[23]), .B(n15344), .C(n10322), .Z(n10343) );
  HS65_LL_NAND2X2 U8371 ( .A(w3[22]), .B(n10343), .Z(n10412) );
  HS65_LL_NAND2AX4 U8372 ( .A(n7733), .B(n7752), .Z(n15045) );
  HS65_LL_NOR2X2 U8373 ( .A(w3[23]), .B(n15045), .Z(n8033) );
  HS65_LL_NOR3X1 U8374 ( .A(w3[17]), .B(w3[22]), .C(n15691), .Z(n7764) );
  HS65_LL_IVX2 U8375 ( .A(n7764), .Z(n7747) );
  HS65_LL_NOR2X2 U8376 ( .A(n7734), .B(n7747), .Z(n7749) );
  HS65_LL_NOR2X2 U8377 ( .A(n15048), .B(n10322), .Z(n10490) );
  HS65_LL_NAND2X2 U8378 ( .A(n10422), .B(n7735), .Z(n10341) );
  HS65_LL_NAND2X2 U8379 ( .A(n7751), .B(n8026), .Z(n8024) );
  HS65_LL_NAND2X2 U8380 ( .A(n10341), .B(n8024), .Z(n10407) );
  HS65_LL_IVX2 U8381 ( .A(n10407), .Z(n15075) );
  HS65_LL_NAND2X2 U8382 ( .A(n7751), .B(n7753), .Z(n10494) );
  HS65_LL_NAND4ABX3 U8383 ( .A(n7749), .B(n10490), .C(n15075), .D(n10494), .Z(
        n7736) );
  HS65_LL_NOR4ABX2 U8384 ( .A(n10442), .B(n10412), .C(n8033), .D(n7736), .Z(
        n10478) );
  HS65_LL_IVX2 U8385 ( .A(n15046), .Z(n8022) );
  HS65_LL_NAND2X2 U8386 ( .A(n8022), .B(n7764), .Z(n10516) );
  HS65_LL_IVX2 U8387 ( .A(n10516), .Z(n10375) );
  HS65_LL_IVX2 U8388 ( .A(n7761), .Z(n7743) );
  HS65_LL_NAND3X2 U8389 ( .A(n15691), .B(n10324), .C(n7743), .Z(n8028) );
  HS65_LL_IVX2 U8390 ( .A(n8028), .Z(n8032) );
  HS65_LL_NAND3X2 U8391 ( .A(w3[17]), .B(n10422), .C(n15691), .Z(n8013) );
  HS65_LL_NOR2X2 U8392 ( .A(n8018), .B(n7747), .Z(n15058) );
  HS65_LL_IVX2 U8393 ( .A(n15058), .Z(n8003) );
  HS65_LL_NAND2X2 U8394 ( .A(n7737), .B(n8022), .Z(n10486) );
  HS65_LL_NAND3X2 U8395 ( .A(n8013), .B(n8003), .C(n10486), .Z(n10467) );
  HS65_LL_NOR3X1 U8396 ( .A(n10375), .B(n8032), .C(n10467), .Z(n10398) );
  HS65_LL_NAND3X2 U8397 ( .A(n10414), .B(n10478), .C(n10398), .Z(n7771) );
  HS65_LL_NOR2X2 U8398 ( .A(w3[18]), .B(w3[20]), .Z(n15088) );
  HS65_LL_IVX2 U8399 ( .A(n8026), .Z(n8005) );
  HS65_LL_NOR2X2 U8400 ( .A(n8005), .B(n10524), .Z(n10321) );
  HS65_LL_IVX2 U8401 ( .A(n7763), .Z(n8006) );
  HS65_LL_NOR3X1 U8402 ( .A(w3[21]), .B(n8006), .C(n8005), .Z(n10449) );
  HS65_LL_NOR2X2 U8403 ( .A(n7746), .B(n7747), .Z(n10506) );
  HS65_LL_NOR2X2 U8404 ( .A(n10496), .B(n10506), .Z(n7738) );
  HS65_LL_NOR2X2 U8405 ( .A(n8018), .B(n7748), .Z(n10493) );
  HS65_LL_IVX2 U8406 ( .A(n10493), .Z(n10517) );
  HS65_LL_NOR2X2 U8407 ( .A(n10524), .B(n8043), .Z(n10312) );
  HS65_LL_IVX2 U8408 ( .A(n10312), .Z(n8004) );
  HS65_LL_NAND3X2 U8409 ( .A(n7738), .B(n10517), .C(n8004), .Z(n7739) );
  HS65_LL_NOR3X1 U8410 ( .A(n10321), .B(n10449), .C(n7739), .Z(n10431) );
  HS65_LL_NOR2X2 U8411 ( .A(n8035), .B(n7740), .Z(n10469) );
  HS65_LL_NOR3X1 U8412 ( .A(n10340), .B(n10469), .C(n10316), .Z(n8046) );
  HS65_LL_NOR2X2 U8413 ( .A(w3[23]), .B(n8020), .Z(n10511) );
  HS65_LL_NOR3AX2 U8414 ( .A(n8012), .B(n15681), .C(n8005), .Z(n10502) );
  HS65_LL_IVX2 U8415 ( .A(n7751), .Z(n7758) );
  HS65_LL_NOR2X2 U8416 ( .A(n7758), .B(n8043), .Z(n10406) );
  HS65_LL_NOR2X2 U8417 ( .A(n8018), .B(n8005), .Z(n10347) );
  HS65_LL_OR2X4 U8418 ( .A(n10406), .B(n10347), .Z(n10415) );
  HS65_LL_NAND2X2 U8419 ( .A(n7743), .B(n7764), .Z(n10381) );
  HS65_LL_NOR2AX3 U8420 ( .A(n10381), .B(n10484), .Z(n10447) );
  HS65_LL_NOR2X2 U8421 ( .A(n10524), .B(n7740), .Z(n10364) );
  HS65_LL_IVX2 U8422 ( .A(n10364), .Z(n8029) );
  HS65_LL_NOR4ABX2 U8423 ( .A(n10447), .B(n8029), .C(n7749), .D(n10464), .Z(
        n10372) );
  HS65_LL_IVX2 U8424 ( .A(n8024), .Z(n10366) );
  HS65_LL_NOR2X2 U8425 ( .A(n8036), .B(n10322), .Z(n10495) );
  HS65_LL_NAND2X2 U8426 ( .A(w3[21]), .B(n10352), .Z(n10315) );
  HS65_LL_IVX2 U8427 ( .A(n10341), .Z(n8015) );
  HS65_LL_NOR2AX3 U8428 ( .A(n10315), .B(n8015), .Z(n8040) );
  HS65_LL_NAND2X2 U8429 ( .A(n8040), .B(n10486), .Z(n10434) );
  HS65_LL_NOR2X2 U8430 ( .A(n15048), .B(n10524), .Z(n10373) );
  HS65_LL_NOR2X2 U8431 ( .A(n15048), .B(n7761), .Z(n10453) );
  HS65_LL_NOR2X2 U8432 ( .A(n10373), .B(n10453), .Z(n8014) );
  HS65_LL_NAND4ABX3 U8433 ( .A(n10490), .B(n10434), .C(n8028), .D(n8014), .Z(
        n7741) );
  HS65_LL_NOR3X1 U8434 ( .A(n10366), .B(n10495), .C(n7741), .Z(n15072) );
  HS65_LL_NAND4ABX3 U8435 ( .A(n10502), .B(n10415), .C(n10372), .D(n15072), 
        .Z(n7742) );
  HS65_LL_NOR4ABX2 U8436 ( .A(n8046), .B(n10362), .C(n10511), .D(n7742), .Z(
        n7769) );
  HS65_LL_IVX2 U8437 ( .A(w3[18]), .Z(n15785) );
  HS65_LL_NAND2X2 U8438 ( .A(w3[20]), .B(n15785), .Z(n10535) );
  HS65_LL_NAND2X2 U8439 ( .A(w3[18]), .B(w3[20]), .Z(n10527) );
  HS65_LL_IVX2 U8440 ( .A(n10527), .Z(n15086) );
  HS65_LL_NAND2X2 U8441 ( .A(n8022), .B(n7754), .Z(n10361) );
  HS65_LL_IVX2 U8442 ( .A(n10361), .Z(n10468) );
  HS65_LL_NOR2X2 U8443 ( .A(n10459), .B(n10468), .Z(n10455) );
  HS65_LL_NOR2X2 U8444 ( .A(n10524), .B(n7748), .Z(n8038) );
  HS65_LL_AOI12X2 U8445 ( .A(n7743), .B(n10324), .C(n8038), .Z(n10444) );
  HS65_LL_NOR2X2 U8446 ( .A(n8035), .B(n7747), .Z(n15077) );
  HS65_LL_NAND2X2 U8447 ( .A(n7751), .B(n7764), .Z(n15051) );
  HS65_LL_IVX2 U8448 ( .A(n15051), .Z(n10377) );
  HS65_LL_NOR3X1 U8449 ( .A(n15077), .B(n10377), .C(n10490), .Z(n7744) );
  HS65_LL_NAND3X2 U8450 ( .A(n10455), .B(n10444), .C(n7744), .Z(n10533) );
  HS65_LL_IVX2 U8451 ( .A(n10533), .Z(n7745) );
  HS65_LL_OAI21X2 U8452 ( .A(n10523), .B(n7761), .C(n7745), .Z(n8048) );
  HS65_LL_NOR2X2 U8453 ( .A(n8043), .B(n7746), .Z(n10417) );
  HS65_LL_NAND4ABX3 U8454 ( .A(n10373), .B(n10417), .C(n10489), .D(n10486), 
        .Z(n7757) );
  HS65_LL_NOR3X1 U8455 ( .A(w3[21]), .B(n8006), .C(n7747), .Z(n10419) );
  HS65_LL_NOR2X2 U8456 ( .A(n15691), .B(n15045), .Z(n10460) );
  HS65_LL_NOR3X1 U8457 ( .A(n10511), .B(n10419), .C(n10460), .Z(n10487) );
  HS65_LL_NOR2X2 U8458 ( .A(n8018), .B(n8036), .Z(n15062) );
  HS65_LL_NOR2X2 U8459 ( .A(n15062), .B(n10321), .Z(n7750) );
  HS65_LL_NOR2X2 U8460 ( .A(n8035), .B(n7748), .Z(n10320) );
  HS65_LL_NAND2X2 U8461 ( .A(w3[21]), .B(n7749), .Z(n8027) );
  HS65_LL_IVX2 U8462 ( .A(n8027), .Z(n10326) );
  HS65_LL_NOR4ABX2 U8463 ( .A(n10487), .B(n7750), .C(n10320), .D(n10326), .Z(
        n15069) );
  HS65_LL_NAND2X2 U8464 ( .A(n7751), .B(n8023), .Z(n10522) );
  HS65_LL_IVX2 U8465 ( .A(n10522), .Z(n7759) );
  HS65_LL_NOR2X2 U8466 ( .A(n7759), .B(n10502), .Z(n10368) );
  HS65_LL_NOR2X2 U8467 ( .A(n10443), .B(n10495), .Z(n8045) );
  HS65_LL_NAND3X2 U8468 ( .A(n10368), .B(n8045), .C(n10412), .Z(n10428) );
  HS65_LL_NAND2X2 U8469 ( .A(n7753), .B(n7752), .Z(n8019) );
  HS65_LL_NAND2X2 U8470 ( .A(n10422), .B(n7754), .Z(n10450) );
  HS65_LL_AND2X4 U8471 ( .A(n8019), .B(n10450), .Z(n10504) );
  HS65_LL_NOR2X2 U8472 ( .A(n7758), .B(n15048), .Z(n10365) );
  HS65_LL_AOI12X2 U8473 ( .A(n8022), .B(n8023), .C(n10365), .Z(n10509) );
  HS65_LL_IVX2 U8474 ( .A(n10347), .Z(n7755) );
  HS65_LL_NAND2X2 U8475 ( .A(n7755), .B(n10381), .Z(n10520) );
  HS65_LL_NOR3X1 U8476 ( .A(n10312), .B(n10366), .C(n10520), .Z(n7756) );
  HS65_LL_NAND3X2 U8477 ( .A(n10504), .B(n10509), .C(n7756), .Z(n10331) );
  HS65_LL_NOR2X2 U8478 ( .A(n10428), .B(n10331), .Z(n8042) );
  HS65_LL_NAND4ABX3 U8479 ( .A(n8048), .B(n7757), .C(n15069), .D(n8042), .Z(
        n7767) );
  HS65_LL_NOR2X2 U8480 ( .A(w3[20]), .B(n15785), .Z(n15084) );
  HS65_LL_NOR3X1 U8481 ( .A(w3[23]), .B(n7758), .C(n15344), .Z(n10510) );
  HS65_LL_NAND2X2 U8482 ( .A(w3[22]), .B(n10510), .Z(n10383) );
  HS65_LL_NAND2X2 U8483 ( .A(n15051), .B(n10383), .Z(n8021) );
  HS65_LL_NOR2X2 U8484 ( .A(n8005), .B(n7761), .Z(n15068) );
  HS65_LL_NOR2X2 U8485 ( .A(n10449), .B(n15068), .Z(n8034) );
  HS65_LL_NOR2X2 U8486 ( .A(n15056), .B(n10459), .Z(n10349) );
  HS65_LL_NOR4ABX2 U8487 ( .A(n8034), .B(n10349), .C(n7759), .D(n10484), .Z(
        n7760) );
  HS65_LL_IVX2 U8488 ( .A(n10460), .Z(n10342) );
  HS65_LL_NAND4ABX3 U8489 ( .A(n10415), .B(n8021), .C(n7760), .D(n10342), .Z(
        n10481) );
  HS65_LL_NAND3AX3 U8490 ( .A(n8033), .B(n10446), .C(n10450), .Z(n8011) );
  HS65_LL_NOR2X2 U8491 ( .A(n8036), .B(n7761), .Z(n10374) );
  HS65_LL_NOR2X2 U8492 ( .A(n10322), .B(n7762), .Z(n10492) );
  HS65_LL_IVX2 U8493 ( .A(n10485), .Z(n10367) );
  HS65_LL_AOI12X2 U8494 ( .A(n10422), .B(n8026), .C(n10417), .Z(n10385) );
  HS65_LL_NAND4ABX3 U8495 ( .A(n10374), .B(n10492), .C(n10367), .D(n10385), 
        .Z(n10360) );
  HS65_LL_AOI112X2 U8496 ( .A(n7764), .B(n7763), .C(n10469), .D(n10360), .Z(
        n7765) );
  HS65_LL_NAND4ABX3 U8497 ( .A(n10481), .B(n8011), .C(n15072), .D(n7765), .Z(
        n7766) );
  HS65_LL_AOI22X1 U8498 ( .A(n15086), .B(n7767), .C(n15084), .D(n7766), .Z(
        n7768) );
  HS65_LL_CBI4I1X3 U8499 ( .A(n10431), .B(n7769), .C(n10535), .D(n7768), .Z(
        n7770) );
  HS65_LL_CBI4I6X2 U8500 ( .A(n7772), .B(n7771), .C(n15088), .D(n7770), .Z(
        n7773) );
  HS65_LLS_XOR3X2 U8501 ( .A(w0[25]), .B(n7773), .C(\u0/rcon [25]), .Z(n10084)
         );
  HS65_LL_MUXI21X2 U8502 ( .D0(n15136), .D1(w1[25]), .S0(n10084), .Z(n10403)
         );
  HS65_LL_MUXI21X2 U8503 ( .D0(n15193), .D1(w2[25]), .S0(n10403), .Z(n10546)
         );
  HS65_LL_MUX31X4 U8504 ( .D0(n15250), .D1(w3[25]), .D2(key[25]), .S0(n10546), 
        .S1(n15783), .Z(\u0/N265 ) );
  HS65_LL_IVX2 U8505 ( .A(w1[14]), .Z(n15360) );
  HS65_LL_IVX2 U8506 ( .A(sa23[1]), .Z(n10666) );
  HS65_LL_IVX2 U8507 ( .A(sa23[6]), .Z(n10665) );
  HS65_LL_NOR2X2 U8508 ( .A(n10665), .B(sa23[7]), .Z(n10700) );
  HS65_LL_IVX2 U8509 ( .A(n10700), .Z(n11864) );
  HS65_LL_NOR2X2 U8510 ( .A(n10666), .B(n11864), .Z(n7805) );
  HS65_LL_IVX2 U8511 ( .A(n7805), .Z(n7786) );
  HS65_LL_IVX2 U8512 ( .A(sa23[3]), .Z(n7774) );
  HS65_LL_NOR2X2 U8513 ( .A(sa23[0]), .B(n7774), .Z(n7775) );
  HS65_LL_IVX2 U8514 ( .A(sa23[5]), .Z(n7780) );
  HS65_LL_NAND2X2 U8515 ( .A(n7775), .B(n7780), .Z(n10664) );
  HS65_LL_NOR2X2 U8516 ( .A(n7786), .B(n10664), .Z(n10868) );
  HS65_LL_NAND2X2 U8517 ( .A(sa23[7]), .B(n10665), .Z(n13434) );
  HS65_LL_IVX2 U8518 ( .A(n13434), .Z(n7777) );
  HS65_LL_NAND2X2 U8519 ( .A(sa23[5]), .B(n7775), .Z(n10655) );
  HS65_LL_NOR2X2 U8520 ( .A(sa23[1]), .B(n10655), .Z(n11856) );
  HS65_LL_NAND2X2 U8521 ( .A(n7777), .B(n11856), .Z(n11860) );
  HS65_LL_IVX2 U8522 ( .A(n11860), .Z(n10859) );
  HS65_LL_NOR2X2 U8523 ( .A(n10868), .B(n10859), .Z(n7779) );
  HS65_LL_NOR2X2 U8524 ( .A(sa23[6]), .B(sa23[7]), .Z(n14306) );
  HS65_LL_NAND2X2 U8525 ( .A(sa23[1]), .B(n14306), .Z(n7785) );
  HS65_LL_NAND2X2 U8526 ( .A(sa23[0]), .B(n7774), .Z(n7776) );
  HS65_LL_NOR2X2 U8527 ( .A(sa23[5]), .B(n7776), .Z(n7801) );
  HS65_LL_IVX2 U8528 ( .A(n7801), .Z(n13435) );
  HS65_LL_NOR2X2 U8529 ( .A(n7785), .B(n13435), .Z(n12213) );
  HS65_LL_NAND3X2 U8530 ( .A(sa23[1]), .B(sa23[6]), .C(sa23[7]), .Z(n10690) );
  HS65_LL_NOR2X2 U8531 ( .A(n10690), .B(n10655), .Z(n13446) );
  HS65_LL_NOR3X1 U8532 ( .A(sa23[1]), .B(sa23[6]), .C(sa23[7]), .Z(n10696) );
  HS65_LL_NAND2X2 U8533 ( .A(n7775), .B(n10696), .Z(n7783) );
  HS65_LL_NOR2X2 U8534 ( .A(sa23[5]), .B(n7783), .Z(n13433) );
  HS65_LL_NOR3X1 U8535 ( .A(n12213), .B(n13446), .C(n13433), .Z(n7778) );
  HS65_LL_IVX2 U8536 ( .A(n7776), .Z(n10874) );
  HS65_LL_NAND2X2 U8537 ( .A(sa23[5]), .B(n10874), .Z(n10842) );
  HS65_LL_NAND2X2 U8538 ( .A(sa23[1]), .B(n7777), .Z(n10656) );
  HS65_LL_NOR2X2 U8539 ( .A(n10842), .B(n10656), .Z(n11827) );
  HS65_LL_IVX2 U8540 ( .A(n11827), .Z(n13447) );
  HS65_LL_NOR3X1 U8541 ( .A(sa23[1]), .B(n10665), .C(n13435), .Z(n12217) );
  HS65_LL_NAND2X2 U8542 ( .A(sa23[7]), .B(n12217), .Z(n12197) );
  HS65_LL_NAND2X2 U8543 ( .A(n13447), .B(n12197), .Z(n14332) );
  HS65_LL_NAND2X2 U8544 ( .A(n7805), .B(n7801), .Z(n11825) );
  HS65_LL_NAND2X2 U8545 ( .A(n10700), .B(n11856), .Z(n11816) );
  HS65_LL_NAND2X2 U8546 ( .A(n11825), .B(n11816), .Z(n12225) );
  HS65_LL_NOR4ABX2 U8547 ( .A(n7779), .B(n7778), .C(n14332), .D(n12225), .Z(
        n14300) );
  HS65_LL_NOR2X2 U8548 ( .A(sa23[3]), .B(sa23[0]), .Z(n10856) );
  HS65_LL_NAND2X2 U8549 ( .A(sa23[5]), .B(n10856), .Z(n11863) );
  HS65_LL_NOR2X2 U8550 ( .A(n7785), .B(n11863), .Z(n10675) );
  HS65_LL_NAND2X2 U8551 ( .A(sa23[3]), .B(sa23[0]), .Z(n14316) );
  HS65_LL_NOR2X2 U8552 ( .A(sa23[5]), .B(n14316), .Z(n7808) );
  HS65_LL_IVX2 U8553 ( .A(n7808), .Z(n7789) );
  HS65_LL_NOR2X2 U8554 ( .A(n7786), .B(n7789), .Z(n13432) );
  HS65_LL_NOR2X2 U8555 ( .A(n7780), .B(n14316), .Z(n10681) );
  HS65_LL_IVX2 U8556 ( .A(n10681), .Z(n7810) );
  HS65_LL_NOR2X2 U8557 ( .A(n7785), .B(n7810), .Z(n12220) );
  HS65_LL_NOR3X1 U8558 ( .A(n10675), .B(n13432), .C(n12220), .Z(n14330) );
  HS65_LL_IVX2 U8559 ( .A(n7785), .Z(n10857) );
  HS65_LL_NAND2X2 U8560 ( .A(n10857), .B(n7808), .Z(n13423) );
  HS65_LL_NOR2X2 U8561 ( .A(n10656), .B(n7810), .Z(n13452) );
  HS65_LL_NOR2X2 U8562 ( .A(n10656), .B(n11863), .Z(n14292) );
  HS65_LL_NOR3AX2 U8563 ( .A(n13423), .B(n13452), .C(n14292), .Z(n10850) );
  HS65_LL_NOR2X2 U8564 ( .A(sa23[1]), .B(n11864), .Z(n12202) );
  HS65_LL_IVX2 U8565 ( .A(n12202), .Z(n14317) );
  HS65_LL_NOR2X2 U8566 ( .A(n7810), .B(n14317), .Z(n10844) );
  HS65_LL_NOR3X1 U8567 ( .A(sa23[5]), .B(sa23[3]), .C(sa23[0]), .Z(n10660) );
  HS65_LL_IVX2 U8568 ( .A(n10660), .Z(n7800) );
  HS65_LL_NAND2X2 U8569 ( .A(sa23[6]), .B(sa23[7]), .Z(n7811) );
  HS65_LL_NOR2X2 U8570 ( .A(sa23[1]), .B(n7811), .Z(n10851) );
  HS65_LL_IVX2 U8571 ( .A(n10851), .Z(n14309) );
  HS65_LL_NOR2X2 U8572 ( .A(n7800), .B(n14309), .Z(n14328) );
  HS65_LL_NOR2X2 U8573 ( .A(n10844), .B(n14328), .Z(n7793) );
  HS65_LL_NAND2X2 U8574 ( .A(n10851), .B(n7808), .Z(n11833) );
  HS65_LL_NAND2X2 U8575 ( .A(n7793), .B(n11833), .Z(n13456) );
  HS65_LL_NOR2X2 U8576 ( .A(n13435), .B(n10690), .Z(n14291) );
  HS65_LL_NOR2X2 U8577 ( .A(sa23[1]), .B(n13434), .Z(n10873) );
  HS65_LL_IVX2 U8578 ( .A(n10873), .Z(n7809) );
  HS65_LL_NOR2X2 U8579 ( .A(n7800), .B(n7809), .Z(n11866) );
  HS65_LL_NOR2X2 U8580 ( .A(n7785), .B(n10664), .Z(n13451) );
  HS65_LL_OR2X4 U8581 ( .A(n11866), .B(n13451), .Z(n11822) );
  HS65_LL_NOR2X2 U8582 ( .A(n10656), .B(n10664), .Z(n13429) );
  HS65_LL_NOR2X2 U8583 ( .A(n10690), .B(n7789), .Z(n13428) );
  HS65_LL_NAND2X2 U8584 ( .A(n10873), .B(n7808), .Z(n10697) );
  HS65_LL_NOR2X2 U8585 ( .A(n10656), .B(n10655), .Z(n11884) );
  HS65_LL_IVX2 U8586 ( .A(n11884), .Z(n14297) );
  HS65_LL_NAND2X2 U8587 ( .A(n10697), .B(n14297), .Z(n7790) );
  HS65_LL_NOR3X1 U8588 ( .A(n13429), .B(n13428), .C(n7790), .Z(n7781) );
  HS65_LL_NAND2X2 U8589 ( .A(n7805), .B(n10681), .Z(n13448) );
  HS65_LL_NAND4ABX3 U8590 ( .A(n14291), .B(n11822), .C(n7781), .D(n13448), .Z(
        n14313) );
  HS65_LL_NOR4ABX2 U8591 ( .A(n14330), .B(n10850), .C(n13456), .D(n14313), .Z(
        n7782) );
  HS65_LL_IVX2 U8592 ( .A(n10690), .Z(n10659) );
  HS65_LL_NAND2X2 U8593 ( .A(n10660), .B(n10659), .Z(n14307) );
  HS65_LL_NOR3X1 U8594 ( .A(sa23[1]), .B(n10665), .C(n10664), .Z(n10667) );
  HS65_LL_NOR2X2 U8595 ( .A(n10842), .B(n14309), .Z(n10691) );
  HS65_LL_NOR2X2 U8596 ( .A(n11863), .B(n7809), .Z(n14299) );
  HS65_LL_NOR2X2 U8597 ( .A(n10691), .B(n14299), .Z(n11891) );
  HS65_LL_NAND3X2 U8598 ( .A(sa23[5]), .B(n10874), .C(n12202), .Z(n14325) );
  HS65_LL_NAND2X2 U8599 ( .A(n11891), .B(n14325), .Z(n10680) );
  HS65_LL_NOR4ABX2 U8600 ( .A(n7782), .B(n14307), .C(n10667), .D(n10680), .Z(
        n7818) );
  HS65_LL_IVX2 U8601 ( .A(sa23[2]), .Z(n7799) );
  HS65_LL_NAND2X2 U8602 ( .A(sa23[4]), .B(n7799), .Z(n11880) );
  HS65_LL_NAND2X2 U8603 ( .A(n12202), .B(n7808), .Z(n10661) );
  HS65_LL_NOR2AX3 U8604 ( .A(n10661), .B(n14292), .Z(n10693) );
  HS65_LL_NOR2X2 U8605 ( .A(n7810), .B(n10690), .Z(n13422) );
  HS65_LL_IVX2 U8606 ( .A(n10842), .Z(n14305) );
  HS65_LL_NAND2X2 U8607 ( .A(n14305), .B(n10857), .Z(n11872) );
  HS65_LL_NAND2X2 U8608 ( .A(n11872), .B(n7783), .Z(n10674) );
  HS65_LL_NOR4ABX2 U8609 ( .A(n10693), .B(n14307), .C(n13422), .D(n10674), .Z(
        n7784) );
  HS65_LL_NAND3AX3 U8610 ( .A(sa23[7]), .B(sa23[1]), .C(n7808), .Z(n10695) );
  HS65_LL_OAI112X1 U8611 ( .A(n7811), .B(n10664), .C(n7784), .D(n10695), .Z(
        n11831) );
  HS65_LL_NAND2X2 U8612 ( .A(n10681), .B(n10696), .Z(n11815) );
  HS65_LL_NAND2X2 U8613 ( .A(n10660), .B(n10696), .Z(n10671) );
  HS65_LL_NAND2X2 U8614 ( .A(n11815), .B(n10671), .Z(n7803) );
  HS65_LL_NAND2X2 U8615 ( .A(n13448), .B(n12197), .Z(n10672) );
  HS65_LL_NOR2X2 U8616 ( .A(n7800), .B(n7785), .Z(n11817) );
  HS65_LL_IVX2 U8617 ( .A(n10656), .Z(n10654) );
  HS65_LL_NAND2X2 U8618 ( .A(n10654), .B(n7801), .Z(n11867) );
  HS65_LL_IVX2 U8619 ( .A(n11867), .Z(n14294) );
  HS65_LL_NOR2X2 U8620 ( .A(n14294), .B(n13429), .Z(n12216) );
  HS65_LL_NOR2X2 U8621 ( .A(n7786), .B(n10842), .Z(n14295) );
  HS65_LL_NOR2X2 U8622 ( .A(n14309), .B(n11863), .Z(n7807) );
  HS65_LL_NOR3X1 U8623 ( .A(n14295), .B(n13452), .C(n7807), .Z(n7787) );
  HS65_LL_NAND3AX3 U8624 ( .A(n11817), .B(n12216), .C(n7787), .Z(n13415) );
  HS65_LL_NAND2X2 U8625 ( .A(n10874), .B(n10696), .Z(n10869) );
  HS65_LL_IVX2 U8626 ( .A(n13451), .Z(n10688) );
  HS65_LL_NAND3X2 U8627 ( .A(sa23[5]), .B(sa23[3]), .C(n10857), .Z(n7802) );
  HS65_LL_NAND3X2 U8628 ( .A(n10869), .B(n10688), .C(n7802), .Z(n7788) );
  HS65_LL_NOR3X1 U8629 ( .A(n13415), .B(n10680), .C(n7788), .Z(n11882) );
  HS65_LL_NOR2X2 U8630 ( .A(n10656), .B(n7789), .Z(n10682) );
  HS65_LL_IVX2 U8631 ( .A(n10696), .Z(n7796) );
  HS65_LL_NOR2X2 U8632 ( .A(n11863), .B(n7796), .Z(n12205) );
  HS65_LL_NOR2X2 U8633 ( .A(n10682), .B(n12205), .Z(n13436) );
  HS65_LL_NAND2X2 U8634 ( .A(n7805), .B(n10856), .Z(n10676) );
  HS65_LL_NOR4ABX2 U8635 ( .A(n13436), .B(n10676), .C(n12213), .D(n7790), .Z(
        n7791) );
  HS65_LL_NOR2X2 U8636 ( .A(n10842), .B(n7809), .Z(n14319) );
  HS65_LL_NOR4ABX2 U8637 ( .A(n11882), .B(n7791), .C(n14291), .D(n14319), .Z(
        n7792) );
  HS65_LL_NAND4ABX3 U8638 ( .A(n7803), .B(n10672), .C(n7793), .D(n7792), .Z(
        n7816) );
  HS65_LL_NOR2X2 U8639 ( .A(sa23[2]), .B(sa23[4]), .Z(n14337) );
  HS65_LL_NOR2X2 U8640 ( .A(sa23[5]), .B(n10869), .Z(n13438) );
  HS65_LL_NOR2X2 U8641 ( .A(sa23[0]), .B(n7802), .Z(n11871) );
  HS65_LL_NAND2X2 U8642 ( .A(n14307), .B(n10671), .Z(n10701) );
  HS65_LL_NAND2X2 U8643 ( .A(n14305), .B(n10696), .Z(n12196) );
  HS65_LL_IVX2 U8644 ( .A(n10664), .Z(n12201) );
  HS65_LL_NAND2X2 U8645 ( .A(n12201), .B(n10873), .Z(n14296) );
  HS65_LL_NAND2X2 U8646 ( .A(n12196), .B(n14296), .Z(n11862) );
  HS65_LL_NOR2X2 U8647 ( .A(n7807), .B(n10682), .Z(n14302) );
  HS65_LL_IVX2 U8648 ( .A(n10844), .Z(n10670) );
  HS65_LL_NAND3AX3 U8649 ( .A(n11862), .B(n14302), .C(n10670), .Z(n7794) );
  HS65_LL_NOR3X1 U8650 ( .A(n11871), .B(n10701), .C(n7794), .Z(n11887) );
  HS65_LL_NOR2X2 U8651 ( .A(n13451), .B(n12205), .Z(n10861) );
  HS65_LL_IVX2 U8652 ( .A(n11863), .Z(n10658) );
  HS65_LL_NAND3X2 U8653 ( .A(sa23[1]), .B(n10700), .C(n10658), .Z(n11845) );
  HS65_LL_NAND3X2 U8654 ( .A(n11887), .B(n10861), .C(n11845), .Z(n7795) );
  HS65_LL_NOR3X1 U8655 ( .A(n13438), .B(n13433), .C(n7795), .Z(n12222) );
  HS65_LL_IVX2 U8656 ( .A(n11825), .Z(n10692) );
  HS65_LL_AOI12X2 U8657 ( .A(n7796), .B(n10690), .C(n10655), .Z(n13441) );
  HS65_LL_NOR3X1 U8658 ( .A(n11817), .B(n10692), .C(n13441), .Z(n10862) );
  HS65_LL_OAI21X2 U8659 ( .A(n10664), .B(n11864), .C(n11833), .Z(n7797) );
  HS65_LL_NOR4ABX2 U8660 ( .A(n10862), .B(n10850), .C(n10672), .D(n7797), .Z(
        n7798) );
  HS65_LL_NOR2X2 U8661 ( .A(n13435), .B(n14317), .Z(n10687) );
  HS65_LL_IVX2 U8662 ( .A(n10675), .Z(n12206) );
  HS65_LL_NAND2X2 U8663 ( .A(n10661), .B(n12206), .Z(n11843) );
  HS65_LL_NOR4ABX2 U8664 ( .A(n7798), .B(n14297), .C(n10687), .D(n11843), .Z(
        n7814) );
  HS65_LL_NOR2X2 U8665 ( .A(n7799), .B(sa23[4]), .Z(n14333) );
  HS65_LL_IVX2 U8666 ( .A(n14333), .Z(n12229) );
  HS65_LL_AOI12X2 U8667 ( .A(n11864), .B(n7809), .C(n7800), .Z(n10871) );
  HS65_LL_NAND2X2 U8668 ( .A(n7801), .B(n10873), .Z(n11875) );
  HS65_LL_NAND4ABX3 U8669 ( .A(n11827), .B(n10871), .C(n11845), .D(n11875), 
        .Z(n13427) );
  HS65_LL_IVX2 U8670 ( .A(n7802), .Z(n7804) );
  HS65_LL_AOI112X2 U8671 ( .A(n11856), .B(n10665), .C(n7804), .D(n7803), .Z(
        n7806) );
  HS65_LL_IVX2 U8672 ( .A(n10655), .Z(n10852) );
  HS65_LL_NAND2X2 U8673 ( .A(n7805), .B(n10852), .Z(n11841) );
  HS65_LL_NAND4ABX3 U8674 ( .A(n10691), .B(n13427), .C(n7806), .D(n11841), .Z(
        n12209) );
  HS65_LL_NOR2X2 U8675 ( .A(n10842), .B(n10690), .Z(n12200) );
  HS65_LL_NOR2X2 U8676 ( .A(n12200), .B(n10844), .Z(n11819) );
  HS65_LL_NOR2X2 U8677 ( .A(n7807), .B(n10687), .Z(n10678) );
  HS65_LL_NAND3X2 U8678 ( .A(n11819), .B(n10678), .C(n14297), .Z(n13444) );
  HS65_LL_NAND2X2 U8679 ( .A(n10696), .B(n7808), .Z(n11844) );
  HS65_LL_NAND2X2 U8680 ( .A(n11844), .B(n14307), .Z(n11854) );
  HS65_LL_NOR2X2 U8681 ( .A(n7810), .B(n7809), .Z(n11818) );
  HS65_LL_IVX2 U8682 ( .A(n11818), .Z(n10698) );
  HS65_LL_OAI21X2 U8683 ( .A(n7811), .B(n10655), .C(n10698), .Z(n11870) );
  HS65_LL_NOR2X2 U8684 ( .A(n14295), .B(n12213), .Z(n10689) );
  HS65_LL_NAND4ABX3 U8685 ( .A(n11854), .B(n11870), .C(n10689), .D(n10688), 
        .Z(n7812) );
  HS65_LL_NAND2X2 U8686 ( .A(sa23[2]), .B(sa23[4]), .Z(n11888) );
  HS65_LL_IVX2 U8687 ( .A(n11888), .Z(n14335) );
  HS65_LL_OAI13X1 U8688 ( .A(n12209), .B(n13444), .C(n7812), .D(n14335), .Z(
        n7813) );
  HS65_LL_CBI4I1X3 U8689 ( .A(n12222), .B(n7814), .C(n12229), .D(n7813), .Z(
        n7815) );
  HS65_LL_CBI4I6X2 U8690 ( .A(n11831), .B(n7816), .C(n14337), .D(n7815), .Z(
        n7817) );
  HS65_LL_CBI4I1X3 U8691 ( .A(n14300), .B(n7818), .C(n11880), .D(n7817), .Z(
        n14983) );
  HS65_LL_IVX2 U8692 ( .A(n14983), .Z(n15361) );
  HS65_LL_IVX2 U8693 ( .A(sa30[0]), .Z(n7819) );
  HS65_LL_NOR2X2 U8694 ( .A(n7819), .B(sa30[5]), .Z(n7820) );
  HS65_LL_IVX2 U8695 ( .A(n7820), .Z(n10146) );
  HS65_LL_NAND3X2 U8696 ( .A(sa30[6]), .B(sa30[7]), .C(sa30[1]), .Z(n10171) );
  HS65_LL_IVX2 U8697 ( .A(sa30[6]), .Z(n7830) );
  HS65_LL_IVX2 U8698 ( .A(sa30[7]), .Z(n10907) );
  HS65_LL_NAND2X2 U8699 ( .A(sa30[1]), .B(n10907), .Z(n12844) );
  HS65_LL_NOR2X2 U8700 ( .A(n7830), .B(n12844), .Z(n7839) );
  HS65_LL_NAND3X2 U8701 ( .A(sa30[3]), .B(sa30[5]), .C(n7839), .Z(n14652) );
  HS65_LL_NOR2X2 U8702 ( .A(n7819), .B(n14652), .Z(n7905) );
  HS65_LL_NAND2X2 U8703 ( .A(n7819), .B(sa30[5]), .Z(n7823) );
  HS65_LL_IVX2 U8704 ( .A(n7823), .Z(n10143) );
  HS65_LL_NAND2X2 U8705 ( .A(sa30[3]), .B(n10143), .Z(n7917) );
  HS65_LL_IVX2 U8706 ( .A(sa30[1]), .Z(n7906) );
  HS65_LL_NAND2X2 U8707 ( .A(sa30[7]), .B(n7830), .Z(n7845) );
  HS65_LL_NOR2X2 U8708 ( .A(n7906), .B(n7845), .Z(n7915) );
  HS65_LL_IVX2 U8709 ( .A(n7915), .Z(n10145) );
  HS65_LL_NOR2X2 U8710 ( .A(n7917), .B(n10145), .Z(n11124) );
  HS65_LL_NOR2X2 U8711 ( .A(n7905), .B(n11124), .Z(n7828) );
  HS65_LL_NOR3X1 U8712 ( .A(sa30[3]), .B(sa30[5]), .C(sa30[0]), .Z(n7916) );
  HS65_LL_IVX2 U8713 ( .A(n7845), .Z(n14658) );
  HS65_LL_NAND2X2 U8714 ( .A(n14658), .B(n7906), .Z(n7837) );
  HS65_LL_IVX2 U8715 ( .A(n7837), .Z(n7943) );
  HS65_LL_NAND2X2 U8716 ( .A(n7916), .B(n7943), .Z(n12812) );
  HS65_LL_NAND2X2 U8717 ( .A(sa30[3]), .B(n7820), .Z(n10155) );
  HS65_LL_NOR2X2 U8718 ( .A(n10155), .B(n7837), .Z(n7935) );
  HS65_LL_NOR2X2 U8719 ( .A(sa30[5]), .B(sa30[0]), .Z(n7821) );
  HS65_LL_NAND2X2 U8720 ( .A(sa30[3]), .B(n7821), .Z(n7848) );
  HS65_LL_NOR2X2 U8721 ( .A(n7848), .B(n10145), .Z(n12826) );
  HS65_LL_IVX2 U8722 ( .A(n12826), .Z(n12172) );
  HS65_LL_IVX2 U8723 ( .A(n7848), .Z(n7851) );
  HS65_LL_NOR2X2 U8724 ( .A(sa30[6]), .B(n12844), .Z(n7903) );
  HS65_LL_NAND2X2 U8725 ( .A(n7851), .B(n7903), .Z(n10894) );
  HS65_LL_NAND2X2 U8726 ( .A(n12172), .B(n10894), .Z(n14648) );
  HS65_LL_NOR4ABX2 U8727 ( .A(n7828), .B(n12812), .C(n7935), .D(n14648), .Z(
        n7822) );
  HS65_LL_OAI21X2 U8728 ( .A(n10146), .B(n10171), .C(n7822), .Z(n10886) );
  HS65_LL_IVX2 U8729 ( .A(sa30[3]), .Z(n10163) );
  HS65_LL_NAND2X2 U8730 ( .A(sa30[5]), .B(sa30[0]), .Z(n12150) );
  HS65_LL_NOR2X2 U8731 ( .A(n10163), .B(n12150), .Z(n10158) );
  HS65_LL_IVX2 U8732 ( .A(n10155), .Z(n12843) );
  HS65_LL_NAND2X2 U8733 ( .A(n12843), .B(n7903), .Z(n10901) );
  HS65_LL_IVX2 U8734 ( .A(n10901), .Z(n14681) );
  HS65_LL_AOI12X2 U8735 ( .A(n7915), .B(n10158), .C(n14681), .Z(n7923) );
  HS65_LL_NOR2X2 U8736 ( .A(sa30[3]), .B(n7823), .Z(n14659) );
  HS65_LL_NAND3X2 U8737 ( .A(sa30[1]), .B(n14658), .C(n14659), .Z(n12184) );
  HS65_LL_NAND2X2 U8738 ( .A(n7923), .B(n12184), .Z(n10921) );
  HS65_LL_NAND2X2 U8739 ( .A(sa30[6]), .B(n7906), .Z(n7824) );
  HS65_LL_IVX2 U8740 ( .A(n7824), .Z(n10159) );
  HS65_LL_NAND2X2 U8741 ( .A(n7851), .B(n10159), .Z(n7930) );
  HS65_LL_IVX2 U8742 ( .A(n7930), .Z(n7827) );
  HS65_LL_NAND2X2 U8743 ( .A(n14659), .B(n7903), .Z(n10895) );
  HS65_LL_NAND2X2 U8744 ( .A(n7903), .B(n10158), .Z(n7941) );
  HS65_LL_NAND2X2 U8745 ( .A(n12843), .B(n7839), .Z(n12173) );
  HS65_LL_NAND3X2 U8746 ( .A(n10895), .B(n7941), .C(n12173), .Z(n12819) );
  HS65_LL_IVX2 U8747 ( .A(n10171), .Z(n7849) );
  HS65_LL_NAND2X2 U8748 ( .A(n7916), .B(n7849), .Z(n7909) );
  HS65_LL_NOR2X2 U8749 ( .A(sa30[7]), .B(n7824), .Z(n7919) );
  HS65_LL_NOR2X2 U8750 ( .A(sa30[3]), .B(n12150), .Z(n7847) );
  HS65_LL_NAND2X2 U8751 ( .A(n7919), .B(n7847), .Z(n10909) );
  HS65_LL_IVX2 U8752 ( .A(n10909), .Z(n14674) );
  HS65_LL_NAND2X2 U8753 ( .A(sa30[6]), .B(sa30[7]), .Z(n12842) );
  HS65_LL_NOR2X2 U8754 ( .A(sa30[1]), .B(n12842), .Z(n12166) );
  HS65_LL_NAND2X2 U8755 ( .A(n12166), .B(n7847), .Z(n10883) );
  HS65_LL_NAND2X2 U8756 ( .A(n14659), .B(n7943), .Z(n10916) );
  HS65_LL_NAND2X2 U8757 ( .A(n10883), .B(n10916), .Z(n12831) );
  HS65_LL_NOR2X2 U8758 ( .A(n14674), .B(n12831), .Z(n7928) );
  HS65_LL_NAND4ABX3 U8759 ( .A(n7827), .B(n12819), .C(n7909), .D(n7928), .Z(
        n7826) );
  HS65_LL_IVX2 U8760 ( .A(n7839), .Z(n7836) );
  HS65_LL_NOR2X2 U8761 ( .A(sa30[3]), .B(n10146), .Z(n12167) );
  HS65_LL_IVX2 U8762 ( .A(n12167), .Z(n7838) );
  HS65_LL_NOR2X2 U8763 ( .A(n7836), .B(n7838), .Z(n11117) );
  HS65_LL_IVX2 U8764 ( .A(n12166), .Z(n7918) );
  HS65_LL_NOR2X2 U8765 ( .A(n7918), .B(n7838), .Z(n12176) );
  HS65_LL_NOR2X2 U8766 ( .A(n7917), .B(n10171), .Z(n14649) );
  HS65_LL_NOR3X1 U8767 ( .A(n11117), .B(n12176), .C(n14649), .Z(n7829) );
  HS65_LL_IVX2 U8768 ( .A(n7917), .Z(n12168) );
  HS65_LL_NAND2X2 U8769 ( .A(n12168), .B(n7943), .Z(n10906) );
  HS65_LL_NOR2X2 U8770 ( .A(n7848), .B(n7836), .Z(n11125) );
  HS65_LL_NAND3X2 U8771 ( .A(n7830), .B(n10907), .C(n7906), .Z(n7920) );
  HS65_LL_IVX2 U8772 ( .A(n7920), .Z(n10164) );
  HS65_LL_NAND2X2 U8773 ( .A(n7851), .B(n10164), .Z(n11118) );
  HS65_LL_IVX2 U8774 ( .A(n11118), .Z(n14661) );
  HS65_LL_NAND2X2 U8775 ( .A(n7847), .B(n7915), .Z(n7841) );
  HS65_LL_IVX2 U8776 ( .A(n7841), .Z(n12834) );
  HS65_LL_NOR2X2 U8777 ( .A(n14661), .B(n12834), .Z(n7922) );
  HS65_LL_NAND2X2 U8778 ( .A(n7903), .B(n12167), .Z(n7914) );
  HS65_LL_NAND2X2 U8779 ( .A(n7919), .B(n12168), .Z(n12811) );
  HS65_LL_NAND3X2 U8780 ( .A(n7922), .B(n7914), .C(n12811), .Z(n7825) );
  HS65_LL_NOR4ABX2 U8781 ( .A(n7829), .B(n10906), .C(n11125), .D(n7825), .Z(
        n14673) );
  HS65_LL_NAND2X2 U8782 ( .A(n12843), .B(n12166), .Z(n12178) );
  HS65_LL_NAND2X2 U8783 ( .A(n7919), .B(n10158), .Z(n12177) );
  HS65_LL_IVX2 U8784 ( .A(n12177), .Z(n10920) );
  HS65_LL_NAND2X2 U8785 ( .A(n12166), .B(n7916), .Z(n7846) );
  HS65_LL_IVX2 U8786 ( .A(n7846), .Z(n12156) );
  HS65_LL_NOR3AX2 U8787 ( .A(n12178), .B(n10920), .C(n12156), .Z(n14650) );
  HS65_LL_NAND4ABX3 U8788 ( .A(n10921), .B(n7826), .C(n14673), .D(n14650), .Z(
        n7861) );
  HS65_LL_IVX2 U8789 ( .A(sa30[4]), .Z(n7834) );
  HS65_LL_NOR2X2 U8790 ( .A(sa30[2]), .B(n7834), .Z(n14685) );
  HS65_LL_IVX2 U8791 ( .A(n10895), .Z(n12832) );
  HS65_LL_AOI112X2 U8792 ( .A(n12843), .B(n10159), .C(n12832), .D(n10921), .Z(
        n7833) );
  HS65_LL_NAND2X2 U8793 ( .A(n7919), .B(n12167), .Z(n12174) );
  HS65_LL_NAND2X2 U8794 ( .A(n7827), .B(n10907), .Z(n12161) );
  HS65_LL_IVX2 U8795 ( .A(n12161), .Z(n7901) );
  HS65_LL_NOR4ABX2 U8796 ( .A(n7828), .B(n12174), .C(n11125), .D(n7901), .Z(
        n7832) );
  HS65_LL_NAND2X2 U8797 ( .A(n10164), .B(n12168), .Z(n12851) );
  HS65_LL_NAND2X2 U8798 ( .A(n7903), .B(n7916), .Z(n10153) );
  HS65_LL_NAND3X2 U8799 ( .A(n7829), .B(n12851), .C(n10153), .Z(n12823) );
  HS65_LL_NAND2X2 U8800 ( .A(n10164), .B(n12167), .Z(n10889) );
  HS65_LL_NAND2X2 U8801 ( .A(n10889), .B(n10894), .Z(n7854) );
  HS65_LL_IVX2 U8802 ( .A(n14659), .Z(n10908) );
  HS65_LL_NOR3X1 U8803 ( .A(n7830), .B(n12844), .C(n10908), .Z(n7936) );
  HS65_LL_IVX2 U8804 ( .A(n7936), .Z(n7840) );
  HS65_LL_OAI21X2 U8805 ( .A(n10908), .B(n7920), .C(n7840), .Z(n11127) );
  HS65_LL_NAND3X2 U8806 ( .A(sa30[3]), .B(sa30[5]), .C(n7903), .Z(n7852) );
  HS65_LL_NOR2X2 U8807 ( .A(sa30[0]), .B(n7852), .Z(n11129) );
  HS65_LL_NAND2X2 U8808 ( .A(n12166), .B(n14659), .Z(n7926) );
  HS65_LL_NAND2X2 U8809 ( .A(n12843), .B(n7915), .Z(n10902) );
  HS65_LL_NAND2X2 U8810 ( .A(n7926), .B(n10902), .Z(n12813) );
  HS65_LL_NAND2X2 U8811 ( .A(n10164), .B(n7847), .Z(n12169) );
  HS65_LL_NAND2X2 U8812 ( .A(n7851), .B(n7943), .Z(n7933) );
  HS65_LL_NAND2X2 U8813 ( .A(n12169), .B(n7933), .Z(n10152) );
  HS65_LL_NAND2X2 U8814 ( .A(n10164), .B(n7916), .Z(n7912) );
  HS65_LL_NAND4ABX3 U8815 ( .A(n10920), .B(n10152), .C(n7909), .D(n7912), .Z(
        n7831) );
  HS65_LL_NOR3X1 U8816 ( .A(n11129), .B(n12813), .C(n7831), .Z(n11112) );
  HS65_LL_NAND4ABX3 U8817 ( .A(n7854), .B(n11127), .C(n11112), .D(n11118), .Z(
        n12153) );
  HS65_LL_NOR4ABX2 U8818 ( .A(n7833), .B(n7832), .C(n12823), .D(n12153), .Z(
        n7859) );
  HS65_LL_NAND2X2 U8819 ( .A(sa30[2]), .B(n7834), .Z(n12849) );
  HS65_LL_NAND2X2 U8820 ( .A(n12174), .B(n7926), .Z(n7835) );
  HS65_LL_NAND2X2 U8821 ( .A(n7847), .B(n7849), .Z(n12830) );
  HS65_LL_NAND4ABX3 U8822 ( .A(n11124), .B(n7835), .C(n12177), .D(n12830), .Z(
        n14660) );
  HS65_LL_OA12X4 U8823 ( .A(n10155), .B(n7920), .C(n7909), .Z(n10157) );
  HS65_LL_NAND2X2 U8824 ( .A(n10158), .B(n7943), .Z(n10882) );
  HS65_LL_NAND2X2 U8825 ( .A(n10157), .B(n10882), .Z(n10165) );
  HS65_LL_NOR2X2 U8826 ( .A(n7917), .B(n12842), .Z(n11131) );
  HS65_LL_NAND2X2 U8827 ( .A(n7847), .B(n7839), .Z(n10917) );
  HS65_LL_NAND2X2 U8828 ( .A(n10917), .B(n7914), .Z(n7904) );
  HS65_LL_NAND2X2 U8829 ( .A(n10164), .B(n10158), .Z(n10915) );
  HS65_LL_NAND2X2 U8830 ( .A(n10883), .B(n10915), .Z(n7843) );
  HS65_LL_NOR2X2 U8831 ( .A(n7917), .B(n7836), .Z(n12846) );
  HS65_LL_NAND2X2 U8832 ( .A(n7919), .B(n7916), .Z(n12829) );
  HS65_LL_NOR2X2 U8833 ( .A(n7838), .B(n7837), .Z(n10900) );
  HS65_LL_IVX2 U8834 ( .A(n10900), .Z(n10147) );
  HS65_LL_NAND2X2 U8835 ( .A(n12829), .B(n10147), .Z(n12841) );
  HS65_LL_NAND2X2 U8836 ( .A(n7916), .B(n7839), .Z(n12827) );
  HS65_LL_NAND2X2 U8837 ( .A(n12827), .B(n12812), .Z(n10890) );
  HS65_LL_NAND4ABX3 U8838 ( .A(n12841), .B(n10890), .C(n7841), .D(n7840), .Z(
        n14680) );
  HS65_LL_NAND4ABX3 U8839 ( .A(n12846), .B(n14680), .C(n10906), .D(n7912), .Z(
        n7842) );
  HS65_LL_NOR4ABX2 U8840 ( .A(n12851), .B(n7852), .C(n7843), .D(n7842), .Z(
        n12158) );
  HS65_LL_NAND4ABX3 U8841 ( .A(n11131), .B(n7904), .C(n12158), .D(n10894), .Z(
        n7844) );
  HS65_LL_NAND2X2 U8842 ( .A(sa30[4]), .B(sa30[2]), .Z(n14687) );
  HS65_LL_IVX2 U8843 ( .A(n14687), .Z(n12192) );
  HS65_LL_OAI13X1 U8844 ( .A(n14660), .B(n10165), .C(n7844), .D(n12192), .Z(
        n7858) );
  HS65_LL_AND2X4 U8845 ( .A(n7847), .B(n7943), .Z(n10154) );
  HS65_LL_NOR2X2 U8846 ( .A(n10154), .B(n11127), .Z(n10904) );
  HS65_LL_OAI112X1 U8847 ( .A(n7845), .B(n10155), .C(n10904), .D(n12827), .Z(
        n7856) );
  HS65_LL_NAND3X2 U8848 ( .A(n7914), .B(n10915), .C(n7846), .Z(n12182) );
  HS65_LL_NAND2X2 U8849 ( .A(n7919), .B(n12843), .Z(n7913) );
  HS65_LL_NAND2X2 U8850 ( .A(n11118), .B(n7913), .Z(n10161) );
  HS65_LL_NOR2X2 U8851 ( .A(n10155), .B(n12844), .Z(n14665) );
  HS65_LL_NAND2X2 U8852 ( .A(n7847), .B(n7903), .Z(n10923) );
  HS65_LL_NAND2X2 U8853 ( .A(n10923), .B(n7909), .Z(n10149) );
  HS65_LL_NOR2X2 U8854 ( .A(n7848), .B(n10171), .Z(n14655) );
  HS65_LL_NAND2X2 U8855 ( .A(n7849), .B(n10158), .Z(n12149) );
  HS65_LL_IVX2 U8856 ( .A(n12149), .Z(n14675) );
  HS65_LL_NOR2X2 U8857 ( .A(n14655), .B(n14675), .Z(n10898) );
  HS65_LL_NAND4ABX3 U8858 ( .A(n14665), .B(n10149), .C(n10898), .D(n12184), 
        .Z(n7850) );
  HS65_LL_NAND2X2 U8859 ( .A(n7851), .B(n12166), .Z(n7939) );
  HS65_LL_NAND4ABX3 U8860 ( .A(n10161), .B(n7850), .C(n7939), .D(n12851), .Z(
        n12855) );
  HS65_LL_NAND4ABX3 U8861 ( .A(n7905), .B(n12176), .C(n12177), .D(n7912), .Z(
        n7934) );
  HS65_LL_NAND2X2 U8862 ( .A(n12167), .B(n7915), .Z(n11126) );
  HS65_LL_NAND2X2 U8863 ( .A(n10917), .B(n11126), .Z(n10167) );
  HS65_LL_OA12X4 U8864 ( .A(n7851), .B(n10158), .C(n7915), .Z(n12160) );
  HS65_LL_NAND4ABX3 U8865 ( .A(n10167), .B(n12160), .C(n10153), .D(n7926), .Z(
        n14670) );
  HS65_LL_NAND3X2 U8866 ( .A(n7928), .B(n12169), .C(n7852), .Z(n7853) );
  HS65_LL_NOR3X1 U8867 ( .A(n14670), .B(n7854), .C(n7853), .Z(n11139) );
  HS65_LL_NOR3X1 U8868 ( .A(n10146), .B(n10171), .C(sa30[3]), .Z(n10168) );
  HS65_LL_NOR2X2 U8869 ( .A(n10168), .B(n11124), .Z(n14676) );
  HS65_LL_NAND4ABX3 U8870 ( .A(n12855), .B(n7934), .C(n11139), .D(n14676), .Z(
        n7855) );
  HS65_LL_NOR2X2 U8871 ( .A(sa30[4]), .B(sa30[2]), .Z(n14683) );
  HS65_LL_OAI13X1 U8872 ( .A(n7856), .B(n12182), .C(n7855), .D(n14683), .Z(
        n7857) );
  HS65_LL_OAI112X1 U8873 ( .A(n7859), .B(n12849), .C(n7858), .D(n7857), .Z(
        n7860) );
  HS65_LL_CBI4I6X2 U8874 ( .A(n10886), .B(n7861), .C(n14685), .D(n7860), .Z(
        n12148) );
  HS65_LL_NAND3X2 U8875 ( .A(sa01[0]), .B(sa01[3]), .C(sa01[5]), .Z(n7888) );
  HS65_LL_IVX2 U8876 ( .A(sa01[6]), .Z(n7862) );
  HS65_LL_IVX2 U8877 ( .A(sa01[1]), .Z(n11773) );
  HS65_LL_NAND3X2 U8878 ( .A(sa01[7]), .B(n7862), .C(n11773), .Z(n10572) );
  HS65_LL_NOR2X2 U8879 ( .A(n7888), .B(n10572), .Z(n10583) );
  HS65_LL_IVX2 U8880 ( .A(sa01[0]), .Z(n7863) );
  HS65_LL_NOR2X2 U8881 ( .A(sa01[3]), .B(n7863), .Z(n10770) );
  HS65_LL_NAND2X2 U8882 ( .A(sa01[5]), .B(n10770), .Z(n10988) );
  HS65_LL_NOR3X1 U8883 ( .A(sa01[6]), .B(n11773), .C(n10988), .Z(n14427) );
  HS65_LL_NAND2X2 U8884 ( .A(sa01[0]), .B(sa01[3]), .Z(n11602) );
  HS65_LL_NOR2X2 U8885 ( .A(sa01[5]), .B(n11602), .Z(n10553) );
  HS65_LL_IVX2 U8886 ( .A(n10572), .Z(n10766) );
  HS65_LL_NAND2X2 U8887 ( .A(n10553), .B(n10766), .Z(n10555) );
  HS65_LL_IVX2 U8888 ( .A(sa01[7]), .Z(n10794) );
  HS65_LL_NAND2X2 U8889 ( .A(sa01[6]), .B(n10794), .Z(n10987) );
  HS65_LL_NOR2X2 U8890 ( .A(sa01[1]), .B(n10987), .Z(n10771) );
  HS65_LL_NAND2X2 U8891 ( .A(n10771), .B(n10553), .Z(n10598) );
  HS65_LL_NOR2X2 U8892 ( .A(sa01[0]), .B(sa01[3]), .Z(n10973) );
  HS65_LL_IVX2 U8893 ( .A(sa01[5]), .Z(n7871) );
  HS65_LL_NAND2X2 U8894 ( .A(n10973), .B(n7871), .Z(n7877) );
  HS65_LL_IVX2 U8895 ( .A(n7877), .Z(n10575) );
  HS65_LL_NOR3X1 U8896 ( .A(sa01[7]), .B(sa01[6]), .C(sa01[1]), .Z(n11077) );
  HS65_LL_NAND2X2 U8897 ( .A(n10575), .B(n11077), .Z(n10787) );
  HS65_LL_NAND2X2 U8898 ( .A(n10598), .B(n10787), .Z(n11007) );
  HS65_LL_NOR2AX3 U8899 ( .A(n10555), .B(n11007), .Z(n10781) );
  HS65_LL_NAND2X2 U8900 ( .A(sa01[5]), .B(n10973), .Z(n10762) );
  HS65_LL_NOR2X2 U8901 ( .A(n11773), .B(n10987), .Z(n10549) );
  HS65_LL_IVX2 U8902 ( .A(n10549), .Z(n7873) );
  HS65_LL_NOR2X2 U8903 ( .A(n10762), .B(n7873), .Z(n10982) );
  HS65_LL_NAND3X2 U8904 ( .A(sa01[7]), .B(sa01[6]), .C(sa01[1]), .Z(n10552) );
  HS65_LL_NAND2X2 U8905 ( .A(n10770), .B(n7871), .Z(n10573) );
  HS65_LL_NOR2X2 U8906 ( .A(n10552), .B(n10573), .Z(n11564) );
  HS65_LL_NAND3X2 U8907 ( .A(sa01[6]), .B(sa01[7]), .C(n11773), .Z(n11601) );
  HS65_LL_NOR2X2 U8908 ( .A(n7877), .B(n11601), .Z(n11581) );
  HS65_LL_NOR3X1 U8909 ( .A(n10982), .B(n11564), .C(n11581), .Z(n10591) );
  HS65_LL_IVX2 U8910 ( .A(n7888), .Z(n7874) );
  HS65_LL_NAND3X2 U8911 ( .A(sa01[7]), .B(sa01[1]), .C(n7862), .Z(n7887) );
  HS65_LL_IVX2 U8912 ( .A(n7887), .Z(n7866) );
  HS65_LL_NAND2X2 U8913 ( .A(n7874), .B(n7866), .Z(n7890) );
  HS65_LL_IVX2 U8914 ( .A(n10573), .Z(n7867) );
  HS65_LL_NAND2X2 U8915 ( .A(n10549), .B(n7867), .Z(n10785) );
  HS65_LL_IVX2 U8916 ( .A(n10785), .Z(n10547) );
  HS65_LL_NAND2X2 U8917 ( .A(n7863), .B(sa01[3]), .Z(n7865) );
  HS65_LL_IVX2 U8918 ( .A(n7865), .Z(n11078) );
  HS65_LL_NAND2X2 U8919 ( .A(n11078), .B(n7871), .Z(n10569) );
  HS65_LL_IVX2 U8920 ( .A(n10569), .Z(n11776) );
  HS65_LL_NAND3X2 U8921 ( .A(sa01[6]), .B(n11776), .C(n11773), .Z(n10558) );
  HS65_LL_NOR2X2 U8922 ( .A(sa01[7]), .B(n10558), .Z(n14437) );
  HS65_LL_NOR4ABX2 U8923 ( .A(n10591), .B(n7890), .C(n10547), .D(n14437), .Z(
        n7864) );
  HS65_LL_NAND4ABX3 U8924 ( .A(n10583), .B(n14427), .C(n10781), .D(n7864), .Z(
        n14415) );
  HS65_LL_IVX2 U8925 ( .A(n11077), .Z(n10567) );
  HS65_LL_NOR2X2 U8926 ( .A(n10988), .B(n10567), .Z(n10999) );
  HS65_LL_IVX2 U8927 ( .A(n10999), .Z(n11071) );
  HS65_LL_NAND2X2 U8928 ( .A(n10575), .B(n10771), .Z(n11004) );
  HS65_LL_NAND2X2 U8929 ( .A(n11071), .B(n11004), .Z(n11804) );
  HS65_LL_NOR2X2 U8930 ( .A(sa01[7]), .B(sa01[6]), .Z(n10566) );
  HS65_LL_NAND2X2 U8931 ( .A(sa01[1]), .B(n10566), .Z(n7891) );
  HS65_LL_NOR2X2 U8932 ( .A(n7891), .B(n10573), .Z(n10589) );
  HS65_LL_NAND2X2 U8933 ( .A(n10575), .B(n10766), .Z(n10763) );
  HS65_LL_NAND2AX4 U8934 ( .A(n10589), .B(n10763), .Z(n7882) );
  HS65_LL_NAND2X2 U8935 ( .A(n7866), .B(n10575), .Z(n11802) );
  HS65_LL_NOR2X2 U8936 ( .A(n7871), .B(n7865), .Z(n11091) );
  HS65_LL_NAND2X2 U8937 ( .A(n7866), .B(n11091), .Z(n14407) );
  HS65_LL_NAND2X2 U8938 ( .A(n11802), .B(n14407), .Z(n11584) );
  HS65_LL_IVX2 U8939 ( .A(n11601), .Z(n7872) );
  HS65_LL_IVX2 U8940 ( .A(n7891), .Z(n10972) );
  HS65_LL_NAND2X2 U8941 ( .A(n10575), .B(n10972), .Z(n11603) );
  HS65_LL_IVX2 U8942 ( .A(n11603), .Z(n11074) );
  HS65_LL_AOI12X2 U8943 ( .A(n11091), .B(n7872), .C(n11074), .Z(n11796) );
  HS65_LL_NAND3X2 U8944 ( .A(n11078), .B(n10766), .C(n7871), .Z(n11583) );
  HS65_LL_NAND4ABX3 U8945 ( .A(n7882), .B(n11584), .C(n11796), .D(n11583), .Z(
        n11576) );
  HS65_LL_NOR2X2 U8946 ( .A(n10762), .B(n10572), .Z(n14416) );
  HS65_LL_IVX2 U8947 ( .A(n14416), .Z(n11586) );
  HS65_LL_NAND2X2 U8948 ( .A(n11091), .B(n10766), .Z(n10580) );
  HS65_LL_IVX2 U8949 ( .A(n10553), .Z(n7878) );
  HS65_LL_NOR2X2 U8950 ( .A(n7878), .B(n10567), .Z(n10985) );
  HS65_LL_NAND2X2 U8951 ( .A(n10771), .B(n7867), .Z(n11094) );
  HS65_LL_IVX2 U8952 ( .A(n11094), .Z(n10778) );
  HS65_LL_NOR2X2 U8953 ( .A(n10569), .B(n11601), .Z(n10595) );
  HS65_LL_NOR2X2 U8954 ( .A(n7887), .B(n10573), .Z(n11597) );
  HS65_LL_NOR2X2 U8955 ( .A(n10595), .B(n11597), .Z(n14412) );
  HS65_LL_IVX2 U8956 ( .A(n10762), .Z(n7868) );
  HS65_LL_NAND2X2 U8957 ( .A(n7868), .B(n10771), .Z(n11780) );
  HS65_LL_NAND4ABX3 U8958 ( .A(n10985), .B(n10778), .C(n14412), .D(n11780), 
        .Z(n11801) );
  HS65_LL_IVX2 U8959 ( .A(n11091), .Z(n14430) );
  HS65_LL_NOR2X2 U8960 ( .A(n7873), .B(n14430), .Z(n11783) );
  HS65_LL_NOR2X2 U8961 ( .A(n10988), .B(n10572), .Z(n11798) );
  HS65_LL_NOR2X2 U8962 ( .A(n11783), .B(n11798), .Z(n10992) );
  HS65_LL_NAND3X2 U8963 ( .A(sa01[3]), .B(sa01[5]), .C(n10566), .Z(n10577) );
  HS65_LL_NOR2X2 U8964 ( .A(n11773), .B(n10577), .Z(n10564) );
  HS65_LL_NAND2X2 U8965 ( .A(sa01[0]), .B(n10564), .Z(n10550) );
  HS65_LL_NAND2X2 U8966 ( .A(n10992), .B(n10550), .Z(n11085) );
  HS65_LL_NOR4ABX2 U8967 ( .A(n11586), .B(n10580), .C(n11801), .D(n11085), .Z(
        n7869) );
  HS65_LL_NAND2X2 U8968 ( .A(sa01[6]), .B(sa01[1]), .Z(n14431) );
  HS65_LL_NOR2X2 U8969 ( .A(n14431), .B(n10569), .Z(n11598) );
  HS65_LL_NAND2X2 U8970 ( .A(sa01[7]), .B(n11598), .Z(n14423) );
  HS65_LL_NAND4ABX3 U8971 ( .A(n11804), .B(n11576), .C(n7869), .D(n14423), .Z(
        n7900) );
  HS65_LL_IVX2 U8972 ( .A(sa01[2]), .Z(n7886) );
  HS65_LL_NAND2X2 U8973 ( .A(sa01[4]), .B(n7886), .Z(n11587) );
  HS65_LL_IVX2 U8974 ( .A(n11587), .Z(n14447) );
  HS65_LL_NOR2X2 U8975 ( .A(n10567), .B(n14430), .Z(n11582) );
  HS65_LL_NAND2AX4 U8976 ( .A(n11582), .B(n10555), .Z(n10981) );
  HS65_LL_NOR2X2 U8977 ( .A(n10569), .B(n7873), .Z(n11790) );
  HS65_LL_NOR2X2 U8978 ( .A(n10583), .B(n11790), .Z(n10768) );
  HS65_LL_NAND3X2 U8979 ( .A(n10768), .B(n10550), .C(n11583), .Z(n7870) );
  HS65_LL_NOR3X1 U8980 ( .A(n14437), .B(n10981), .C(n7870), .Z(n11806) );
  HS65_LL_NOR2X2 U8981 ( .A(n10552), .B(n10762), .Z(n14442) );
  HS65_LL_NOR2X2 U8982 ( .A(n11601), .B(n10988), .Z(n10578) );
  HS65_LL_NOR2X2 U8983 ( .A(n14442), .B(n10578), .Z(n10792) );
  HS65_LL_NOR2X2 U8984 ( .A(n7878), .B(n11601), .Z(n10784) );
  HS65_LL_NAND2X2 U8985 ( .A(n7874), .B(n10771), .Z(n10986) );
  HS65_LL_IVX2 U8986 ( .A(n10986), .Z(n10590) );
  HS65_LL_NOR3X1 U8987 ( .A(n10784), .B(n10590), .C(n11581), .Z(n14432) );
  HS65_LL_NOR2X2 U8988 ( .A(n7887), .B(n10762), .Z(n11573) );
  HS65_LL_IVX2 U8989 ( .A(n10598), .Z(n10563) );
  HS65_LL_NAND3X2 U8990 ( .A(n7871), .B(n10770), .C(n11077), .Z(n7892) );
  HS65_LL_IVX2 U8991 ( .A(n7892), .Z(n11793) );
  HS65_LL_NAND2X2 U8992 ( .A(n7874), .B(n7872), .Z(n10980) );
  HS65_LL_IVX2 U8993 ( .A(n10980), .Z(n10777) );
  HS65_LL_NOR2X2 U8994 ( .A(n7887), .B(n7878), .Z(n10979) );
  HS65_LL_NOR2X2 U8995 ( .A(n10988), .B(n7873), .Z(n10765) );
  HS65_LL_NOR2X2 U8996 ( .A(n10765), .B(n10589), .Z(n10584) );
  HS65_LL_NAND2X2 U8997 ( .A(n7874), .B(n10549), .Z(n10599) );
  HS65_LL_NAND2X2 U8998 ( .A(n10584), .B(n10599), .Z(n10798) );
  HS65_LL_NOR3X1 U8999 ( .A(n10777), .B(n10979), .C(n10798), .Z(n7875) );
  HS65_LL_NAND4ABX3 U9000 ( .A(n10563), .B(n11793), .C(n10785), .D(n7875), .Z(
        n7876) );
  HS65_LL_NOR4ABX2 U9001 ( .A(n10792), .B(n14432), .C(n11573), .D(n7876), .Z(
        n11073) );
  HS65_LL_NOR2X2 U9002 ( .A(n10552), .B(n7877), .Z(n11606) );
  HS65_LL_NOR2X2 U9003 ( .A(sa01[5]), .B(n7891), .Z(n11003) );
  HS65_LL_NOR4ABX2 U9004 ( .A(n10787), .B(n11094), .C(n11606), .D(n11003), .Z(
        n7879) );
  HS65_LL_NOR2X2 U9005 ( .A(n10552), .B(n10988), .Z(n14438) );
  HS65_LL_NOR3X1 U9006 ( .A(sa01[7]), .B(n11773), .C(n7878), .Z(n10596) );
  HS65_LL_NOR2AX3 U9007 ( .A(n10992), .B(n10596), .Z(n14443) );
  HS65_LL_NAND2X2 U9008 ( .A(n14443), .B(n10580), .Z(n11779) );
  HS65_LL_NOR4ABX2 U9009 ( .A(n11073), .B(n7879), .C(n14438), .D(n11779), .Z(
        n7898) );
  HS65_LL_NAND2X2 U9010 ( .A(sa01[2]), .B(sa01[4]), .Z(n11611) );
  HS65_LL_NOR2X2 U9011 ( .A(sa01[2]), .B(sa01[4]), .Z(n14453) );
  HS65_LL_NOR2X2 U9012 ( .A(n7888), .B(n10552), .Z(n10593) );
  HS65_LL_NOR2X2 U9013 ( .A(n10765), .B(n11597), .Z(n11575) );
  HS65_LL_NOR2X2 U9014 ( .A(n10762), .B(n11601), .Z(n10581) );
  HS65_LL_NOR3X1 U9015 ( .A(sa01[6]), .B(n11773), .C(n10569), .Z(n10556) );
  HS65_LL_NAND2X2 U9016 ( .A(sa01[7]), .B(n10556), .Z(n11092) );
  HS65_LL_NAND2X2 U9017 ( .A(n11092), .B(n7890), .Z(n14426) );
  HS65_LL_NOR4ABX2 U9018 ( .A(n11575), .B(n11603), .C(n10581), .D(n14426), .Z(
        n14440) );
  HS65_LL_NOR2X2 U9019 ( .A(n10569), .B(n7891), .Z(n14424) );
  HS65_LL_NOR2X2 U9020 ( .A(n10578), .B(n14416), .Z(n10974) );
  HS65_LL_NAND3X2 U9021 ( .A(sa01[5]), .B(n10771), .C(n10770), .Z(n14411) );
  HS65_LL_NAND2X2 U9022 ( .A(n10974), .B(n14411), .Z(n10559) );
  HS65_LL_NOR3X1 U9023 ( .A(n10564), .B(n14424), .C(n10559), .Z(n7881) );
  HS65_LL_NAND2X2 U9024 ( .A(n10770), .B(n11077), .Z(n7880) );
  HS65_LL_NAND3X2 U9025 ( .A(n14440), .B(n7881), .C(n7880), .Z(n10783) );
  HS65_LL_IVX2 U9026 ( .A(n10784), .Z(n10561) );
  HS65_LL_NAND2X2 U9027 ( .A(n10561), .B(n10580), .Z(n10990) );
  HS65_LL_NAND3X2 U9028 ( .A(n10768), .B(n14423), .C(n11780), .Z(n11096) );
  HS65_LL_NOR3X1 U9029 ( .A(n10990), .B(n11096), .C(n7882), .Z(n7883) );
  HS65_LL_NAND4ABX3 U9030 ( .A(n10593), .B(n10783), .C(n7883), .D(n10558), .Z(
        n11014) );
  HS65_LL_IVX2 U9031 ( .A(n10771), .Z(n11566) );
  HS65_LL_NOR2X2 U9032 ( .A(n11566), .B(n14430), .Z(n11001) );
  HS65_LL_NAND3X2 U9033 ( .A(n10986), .B(n10787), .C(n11583), .Z(n10565) );
  HS65_LL_IVX2 U9034 ( .A(n10565), .Z(n7885) );
  HS65_LL_NOR2X2 U9035 ( .A(n11601), .B(n10573), .Z(n11577) );
  HS65_LL_NOR2AX3 U9036 ( .A(n10599), .B(n11577), .Z(n7884) );
  HS65_LL_NAND4ABX3 U9037 ( .A(n11014), .B(n11001), .C(n7885), .D(n7884), .Z(
        n7896) );
  HS65_LL_NOR2X2 U9038 ( .A(sa01[4]), .B(n7886), .Z(n14449) );
  HS65_LL_NOR2X2 U9039 ( .A(n7887), .B(n10988), .Z(n10574) );
  HS65_LL_IVX2 U9040 ( .A(n10574), .Z(n11579) );
  HS65_LL_NAND2X2 U9041 ( .A(n10575), .B(n10549), .Z(n11792) );
  HS65_LL_NAND2X2 U9042 ( .A(n11579), .B(n11792), .Z(n10991) );
  HS65_LL_NOR2X2 U9043 ( .A(n10988), .B(n7891), .Z(n11805) );
  HS65_LL_AOI12X2 U9044 ( .A(n11078), .B(n11077), .C(n11805), .Z(n10594) );
  HS65_LL_NAND4ABX3 U9045 ( .A(n10985), .B(n10991), .C(n10594), .D(n11780), 
        .Z(n10774) );
  HS65_LL_NOR2X2 U9046 ( .A(n7888), .B(n10567), .Z(n11000) );
  HS65_LL_NOR3X1 U9047 ( .A(n10595), .B(n11000), .C(n10559), .Z(n7889) );
  HS65_LL_IVX2 U9048 ( .A(n10593), .Z(n10786) );
  HS65_LL_NAND2X2 U9049 ( .A(n10786), .B(n10555), .Z(n14446) );
  HS65_LL_NOR4ABX2 U9050 ( .A(n7889), .B(n11094), .C(n10581), .D(n14446), .Z(
        n14433) );
  HS65_LL_NAND2X2 U9051 ( .A(n10553), .B(n10972), .Z(n14408) );
  HS65_LL_NAND2X2 U9052 ( .A(n14408), .B(n7890), .Z(n10551) );
  HS65_LL_OR2X4 U9053 ( .A(n11007), .B(n10777), .Z(n14436) );
  HS65_LL_NOR2X2 U9054 ( .A(n10762), .B(n7891), .Z(n10562) );
  HS65_LL_NOR3X1 U9055 ( .A(n10979), .B(n10562), .C(n11001), .Z(n11089) );
  HS65_LL_IVX2 U9056 ( .A(n11564), .Z(n11574) );
  HS65_LL_NAND3X2 U9057 ( .A(n11089), .B(n7892), .C(n11574), .Z(n7893) );
  HS65_LL_NOR3X1 U9058 ( .A(n10551), .B(n14436), .C(n7893), .Z(n7894) );
  HS65_LL_NAND4ABX3 U9059 ( .A(n11576), .B(n10774), .C(n14433), .D(n7894), .Z(
        n7895) );
  HS65_LL_AOI22X1 U9060 ( .A(n14453), .B(n7896), .C(n14449), .D(n7895), .Z(
        n7897) );
  HS65_LL_CBI4I1X3 U9061 ( .A(n11806), .B(n7898), .C(n11611), .D(n7897), .Z(
        n7899) );
  HS65_LL_CBI4I6X2 U9062 ( .A(n14415), .B(n7900), .C(n14447), .D(n7899), .Z(
        n15125) );
  HS65_LL_NOR2AX3 U9063 ( .A(n7933), .B(n11125), .Z(n10144) );
  HS65_LL_NOR4ABX2 U9064 ( .A(n10144), .B(n7941), .C(n7935), .D(n7901), .Z(
        n7902) );
  HS65_LL_NAND3X2 U9065 ( .A(n7902), .B(n12851), .C(n10882), .Z(n10925) );
  HS65_LL_NAND3X2 U9066 ( .A(n12830), .B(n10906), .C(n7912), .Z(n7911) );
  HS65_LL_NOR2X2 U9067 ( .A(n12846), .B(n10154), .Z(n12821) );
  HS65_LL_NOR2AX3 U9068 ( .A(n12821), .B(n14665), .Z(n11113) );
  HS65_LL_IVX2 U9069 ( .A(n7903), .Z(n12151) );
  HS65_LL_NOR2X2 U9070 ( .A(sa30[5]), .B(n12151), .Z(n12815) );
  HS65_LL_NOR2X2 U9071 ( .A(n7905), .B(n7904), .Z(n11119) );
  HS65_LL_NAND2X2 U9072 ( .A(n12166), .B(n10158), .Z(n12850) );
  HS65_LL_NOR2AX3 U9073 ( .A(n12850), .B(n11117), .Z(n12838) );
  HS65_LL_NAND2X2 U9074 ( .A(n10889), .B(n10902), .Z(n7924) );
  HS65_LL_OAI13X1 U9075 ( .A(n7906), .B(n10907), .C(n10908), .D(n10883), .Z(
        n7907) );
  HS65_LL_NOR4ABX2 U9076 ( .A(n12838), .B(n7913), .C(n7924), .D(n7907), .Z(
        n7908) );
  HS65_LL_NAND3X2 U9077 ( .A(n11119), .B(n14650), .C(n7908), .Z(n12165) );
  HS65_LL_NOR4ABX2 U9078 ( .A(n11113), .B(n7909), .C(n12815), .D(n12165), .Z(
        n7910) );
  HS65_LL_NAND4ABX3 U9079 ( .A(n10925), .B(n7911), .C(n7910), .D(n12174), .Z(
        n7948) );
  HS65_LL_NAND2X2 U9080 ( .A(n7913), .B(n7912), .Z(n14664) );
  HS65_LL_NOR2X2 U9081 ( .A(n10168), .B(n14664), .Z(n10897) );
  HS65_LL_IVX2 U9082 ( .A(n10897), .Z(n7938) );
  HS65_LL_NAND2X2 U9083 ( .A(n7914), .B(n12812), .Z(n7931) );
  HS65_LL_NAND2X2 U9084 ( .A(n7916), .B(n7915), .Z(n12162) );
  HS65_LL_IVX2 U9085 ( .A(n11124), .Z(n10156) );
  HS65_LL_NAND3X2 U9086 ( .A(n12162), .B(n7933), .C(n10156), .Z(n10169) );
  HS65_LL_OAI21X2 U9087 ( .A(n7918), .B(n7917), .C(n10153), .Z(n10893) );
  HS65_LL_NOR3X1 U9088 ( .A(n7931), .B(n10169), .C(n10893), .Z(n10173) );
  HS65_LL_IVX2 U9089 ( .A(n10173), .Z(n7925) );
  HS65_LL_NAND2X2 U9090 ( .A(n7919), .B(n14659), .Z(n12835) );
  HS65_LL_OAI21X2 U9091 ( .A(n10155), .B(n7920), .C(n12835), .Z(n7940) );
  HS65_LL_NAND2X2 U9092 ( .A(n10923), .B(n12827), .Z(n7921) );
  HS65_LL_NOR4ABX2 U9093 ( .A(n7922), .B(n12851), .C(n7940), .D(n7921), .Z(
        n11111) );
  HS65_LL_NAND4ABX3 U9094 ( .A(n7925), .B(n7924), .C(n7923), .D(n11111), .Z(
        n7929) );
  HS65_LL_IVX2 U9095 ( .A(n10915), .Z(n10885) );
  HS65_LL_NOR2X2 U9096 ( .A(n14675), .B(n7935), .Z(n14667) );
  HS65_LL_NAND3X2 U9097 ( .A(n14667), .B(n12174), .C(n7926), .Z(n7927) );
  HS65_LL_NOR4ABX2 U9098 ( .A(n7928), .B(n7939), .C(n10885), .D(n7927), .Z(
        n14651) );
  HS65_LL_NAND2X2 U9099 ( .A(n12850), .B(n12811), .Z(n12180) );
  HS65_LL_NOR2X2 U9100 ( .A(n12832), .B(n12180), .Z(n12157) );
  HS65_LL_NAND4ABX3 U9101 ( .A(n7938), .B(n7929), .C(n14651), .D(n12157), .Z(
        n7947) );
  HS65_LL_IVX2 U9102 ( .A(n12849), .Z(n14691) );
  HS65_LL_NAND2X2 U9103 ( .A(n12835), .B(n10882), .Z(n11128) );
  HS65_LL_NOR3X1 U9104 ( .A(n14655), .B(n11125), .C(n11128), .Z(n12175) );
  HS65_LL_NAND2X2 U9105 ( .A(n12178), .B(n10906), .Z(n12824) );
  HS65_LL_NAND2X2 U9106 ( .A(n12149), .B(n7930), .Z(n10881) );
  HS65_LL_NOR3X1 U9107 ( .A(n12824), .B(n7931), .C(n10881), .Z(n7932) );
  HS65_LL_NAND3X2 U9108 ( .A(n11139), .B(n12175), .C(n7932), .Z(n12845) );
  HS65_LL_NAND4ABX3 U9109 ( .A(n12845), .B(n7934), .C(n7933), .D(n12811), .Z(
        n7946) );
  HS65_LL_OAI112X1 U9110 ( .A(n12150), .B(n10145), .C(n10923), .D(n12161), .Z(
        n14654) );
  HS65_LL_NOR2X2 U9111 ( .A(n11117), .B(n7935), .Z(n12154) );
  HS65_LL_NAND4ABX3 U9112 ( .A(n12156), .B(n7936), .C(n12154), .D(n10882), .Z(
        n7937) );
  HS65_LL_NOR3X1 U9113 ( .A(n7938), .B(n14654), .C(n7937), .Z(n14663) );
  HS65_LL_AND2X4 U9114 ( .A(n7939), .B(n11126), .Z(n14679) );
  HS65_LL_NAND3AX3 U9115 ( .A(n7940), .B(n14679), .C(n12174), .Z(n10899) );
  HS65_LL_NAND2X2 U9116 ( .A(n12829), .B(n12169), .Z(n10922) );
  HS65_LL_NAND4ABX3 U9117 ( .A(n14655), .B(n10922), .C(n12821), .D(n7941), .Z(
        n7942) );
  HS65_LL_AOI112X2 U9118 ( .A(n10143), .B(n7943), .C(n10899), .D(n7942), .Z(
        n7944) );
  HS65_LL_NAND3X2 U9119 ( .A(n10173), .B(n14663), .C(n7944), .Z(n7945) );
  HS65_LL_MX41X4 U9120 ( .D0(n7948), .S0(n12192), .D1(n7947), .S1(n14691), 
        .D2(n7946), .S2(n14683), .D3(n7945), .S3(n14685), .Z(n15445) );
  HS65_LLS_XNOR2X3 U9121 ( .A(n15125), .B(n15445), .Z(n14957) );
  HS65_LL_IVX2 U9122 ( .A(sa12[6]), .Z(n13392) );
  HS65_LL_NOR2X2 U9123 ( .A(sa12[7]), .B(n13392), .Z(n10810) );
  HS65_LL_NAND2X2 U9124 ( .A(sa12[1]), .B(n10810), .Z(n10060) );
  HS65_LL_NOR3X1 U9125 ( .A(sa12[5]), .B(sa12[0]), .C(sa12[3]), .Z(n10956) );
  HS65_LL_IVX2 U9126 ( .A(n10956), .Z(n7988) );
  HS65_LL_NOR2X2 U9127 ( .A(n10060), .B(n7988), .Z(n10829) );
  HS65_LL_IVX2 U9128 ( .A(sa12[0]), .Z(n7949) );
  HS65_LL_NOR2X2 U9129 ( .A(sa12[3]), .B(n7949), .Z(n7974) );
  HS65_LL_NAND2X2 U9130 ( .A(sa12[5]), .B(n7974), .Z(n7959) );
  HS65_LL_NAND3X2 U9131 ( .A(sa12[1]), .B(sa12[7]), .C(n13392), .Z(n7968) );
  HS65_LL_NOR2X2 U9132 ( .A(n7959), .B(n7968), .Z(n10931) );
  HS65_LL_NOR2X2 U9133 ( .A(n10829), .B(n10931), .Z(n10944) );
  HS65_LL_NOR3X1 U9134 ( .A(sa12[1]), .B(sa12[6]), .C(sa12[7]), .Z(n7975) );
  HS65_LL_IVX2 U9135 ( .A(n7975), .Z(n10960) );
  HS65_LL_IVX2 U9136 ( .A(sa12[3]), .Z(n7950) );
  HS65_LL_NOR2X2 U9137 ( .A(n7949), .B(n7950), .Z(n7985) );
  HS65_LL_IVX2 U9138 ( .A(sa12[5]), .Z(n7984) );
  HS65_LL_NAND2X2 U9139 ( .A(n7985), .B(n7984), .Z(n10958) );
  HS65_LL_NOR2X2 U9140 ( .A(n10960), .B(n10958), .Z(n10070) );
  HS65_LL_IVX2 U9141 ( .A(sa12[1]), .Z(n7963) );
  HS65_LL_NAND2X2 U9142 ( .A(n10810), .B(n7963), .Z(n10720) );
  HS65_LL_NOR3X1 U9143 ( .A(sa12[0]), .B(sa12[3]), .C(n7984), .Z(n7967) );
  HS65_LL_IVX2 U9144 ( .A(n7967), .Z(n10051) );
  HS65_LL_NOR2X2 U9145 ( .A(n10720), .B(n10051), .Z(n10930) );
  HS65_LL_NOR2X2 U9146 ( .A(n10070), .B(n10930), .Z(n7990) );
  HS65_LL_NOR2X2 U9147 ( .A(sa12[0]), .B(n7950), .Z(n7951) );
  HS65_LL_NOR3X1 U9148 ( .A(sa12[6]), .B(sa12[7]), .C(n7963), .Z(n7973) );
  HS65_LL_IVX2 U9149 ( .A(n7973), .Z(n10824) );
  HS65_LL_NOR2X2 U9150 ( .A(n10824), .B(n7959), .Z(n10811) );
  HS65_LL_AOI12X2 U9151 ( .A(n7975), .B(n7951), .C(n10811), .Z(n10628) );
  HS65_LL_NAND3X2 U9152 ( .A(n10944), .B(n7990), .C(n10628), .Z(n10723) );
  HS65_LL_NAND2X2 U9153 ( .A(n7975), .B(n10956), .Z(n10614) );
  HS65_LL_IVX2 U9154 ( .A(n10720), .Z(n10957) );
  HS65_LL_IVX2 U9155 ( .A(n10958), .Z(n10741) );
  HS65_LL_NAND2X2 U9156 ( .A(n10957), .B(n10741), .Z(n10963) );
  HS65_LL_NAND2X2 U9157 ( .A(n10614), .B(n10963), .Z(n13377) );
  HS65_LL_IVX2 U9158 ( .A(n10810), .Z(n11024) );
  HS65_LL_NAND2X2 U9159 ( .A(sa12[5]), .B(n7951), .Z(n11025) );
  HS65_LL_NOR3X1 U9160 ( .A(sa12[1]), .B(n11024), .C(n11025), .Z(n11064) );
  HS65_LL_OR2X4 U9161 ( .A(n13377), .B(n11064), .Z(n7953) );
  HS65_LL_IVX2 U9162 ( .A(n7974), .Z(n10719) );
  HS65_LL_NOR2X2 U9163 ( .A(sa12[5]), .B(n10719), .Z(n10052) );
  HS65_LL_NAND2X2 U9164 ( .A(n7973), .B(n10052), .Z(n11022) );
  HS65_LL_NAND2X2 U9165 ( .A(n10956), .B(n7973), .Z(n10948) );
  HS65_LL_NOR2X2 U9166 ( .A(n11025), .B(n7968), .Z(n10638) );
  HS65_LL_IVX2 U9167 ( .A(n10638), .Z(n10725) );
  HS65_LL_NAND3X2 U9168 ( .A(sa12[7]), .B(n7963), .C(n13392), .Z(n7983) );
  HS65_LL_IVX2 U9169 ( .A(n7983), .Z(n10612) );
  HS65_LL_NAND2X2 U9170 ( .A(n10956), .B(n10612), .Z(n7977) );
  HS65_LL_NAND2X2 U9171 ( .A(n10725), .B(n7977), .Z(n10729) );
  HS65_LL_IVX2 U9172 ( .A(n7968), .Z(n7970) );
  HS65_LL_NAND2X2 U9173 ( .A(n10956), .B(n7970), .Z(n11052) );
  HS65_LL_IVX2 U9174 ( .A(n7951), .Z(n7972) );
  HS65_LL_NOR2X2 U9175 ( .A(sa12[5]), .B(n7972), .Z(n10641) );
  HS65_LL_IVX2 U9176 ( .A(n10641), .Z(n10629) );
  HS65_LL_NOR2X2 U9177 ( .A(n10629), .B(n7983), .Z(n7979) );
  HS65_LL_IVX2 U9178 ( .A(n7979), .Z(n10071) );
  HS65_LL_IVX2 U9179 ( .A(sa12[7]), .Z(n10623) );
  HS65_LL_NOR2X2 U9180 ( .A(n10623), .B(n11025), .Z(n10745) );
  HS65_LL_NAND3X2 U9181 ( .A(sa12[6]), .B(n10745), .C(n7963), .Z(n11041) );
  HS65_LL_NAND3X2 U9182 ( .A(n11052), .B(n10071), .C(n11041), .Z(n7952) );
  HS65_LL_NOR4ABX2 U9183 ( .A(n11022), .B(n10948), .C(n10729), .D(n7952), .Z(
        n10065) );
  HS65_LL_NAND2X2 U9184 ( .A(n7975), .B(n10052), .Z(n10806) );
  HS65_LL_NAND4ABX3 U9185 ( .A(n10723), .B(n7953), .C(n10065), .D(n10806), .Z(
        n7999) );
  HS65_LL_NAND2X2 U9186 ( .A(n10957), .B(n10052), .Z(n10637) );
  HS65_LL_NAND2X2 U9187 ( .A(sa12[6]), .B(sa12[7]), .Z(n10630) );
  HS65_LL_NOR2X2 U9188 ( .A(sa12[1]), .B(n10630), .Z(n7989) );
  HS65_LL_NAND2X2 U9189 ( .A(sa12[5]), .B(n7985), .Z(n7969) );
  HS65_LL_NOR2X2 U9190 ( .A(n7969), .B(n10960), .Z(n10951) );
  HS65_LL_NOR2X2 U9191 ( .A(n10958), .B(n7983), .Z(n10716) );
  HS65_LL_OR2X4 U9192 ( .A(n10951), .B(n10716), .Z(n10631) );
  HS65_LL_CBI4I6X2 U9193 ( .A(n7967), .B(n10641), .C(n7989), .D(n10631), .Z(
        n7954) );
  HS65_LL_IVX2 U9194 ( .A(n7959), .Z(n10809) );
  HS65_LL_NAND2X2 U9195 ( .A(n10809), .B(n7989), .Z(n10739) );
  HS65_LL_IVX2 U9196 ( .A(n10739), .Z(n10616) );
  HS65_LL_NOR2X2 U9197 ( .A(n10051), .B(n7983), .Z(n13386) );
  HS65_LL_NOR2X2 U9198 ( .A(n10616), .B(n13386), .Z(n10724) );
  HS65_LL_NAND2X2 U9199 ( .A(n10957), .B(n10809), .Z(n13397) );
  HS65_LL_NAND2X2 U9200 ( .A(n10724), .B(n13397), .Z(n10608) );
  HS65_LL_NOR2X2 U9201 ( .A(n7963), .B(n10630), .Z(n7958) );
  HS65_LL_IVX2 U9202 ( .A(n7958), .Z(n10056) );
  HS65_LL_NOR2X2 U9203 ( .A(n7969), .B(n10056), .Z(n13400) );
  HS65_LL_NOR4ABX2 U9204 ( .A(n10637), .B(n7954), .C(n10608), .D(n13400), .Z(
        n13368) );
  HS65_LL_NAND2X2 U9205 ( .A(sa12[1]), .B(n10741), .Z(n13391) );
  HS65_LL_NOR3X1 U9206 ( .A(sa12[6]), .B(sa12[7]), .C(n13391), .Z(n10711) );
  HS65_LL_NAND3X2 U9207 ( .A(sa12[6]), .B(sa12[7]), .C(n10052), .Z(n10735) );
  HS65_LL_NOR2X2 U9208 ( .A(n7963), .B(n10735), .Z(n10073) );
  HS65_LL_NOR2X2 U9209 ( .A(n10711), .B(n10073), .Z(n13398) );
  HS65_LL_NOR2X2 U9210 ( .A(n10824), .B(n10051), .Z(n10962) );
  HS65_LL_IVX2 U9211 ( .A(n7969), .Z(n7956) );
  HS65_LL_NAND2X2 U9212 ( .A(n7956), .B(n7989), .Z(n7955) );
  HS65_LL_IVX2 U9213 ( .A(n7955), .Z(n10955) );
  HS65_LL_AOI112X2 U9214 ( .A(n7985), .B(n7970), .C(n10962), .D(n10955), .Z(
        n11058) );
  HS65_LL_NAND3X2 U9215 ( .A(n13368), .B(n13398), .C(n11058), .Z(n7998) );
  HS65_LL_IVX2 U9216 ( .A(sa12[4]), .Z(n7991) );
  HS65_LL_NAND2X2 U9217 ( .A(sa12[2]), .B(n7991), .Z(n10750) );
  HS65_LL_IVX2 U9218 ( .A(n10750), .Z(n13410) );
  HS65_LL_NOR2X2 U9219 ( .A(n10051), .B(n7968), .Z(n10606) );
  HS65_LL_IVX2 U9220 ( .A(n10606), .Z(n10822) );
  HS65_LL_NAND2X2 U9221 ( .A(n10963), .B(n10822), .Z(n10624) );
  HS65_LL_NAND2X2 U9222 ( .A(n10741), .B(n7970), .Z(n11030) );
  HS65_LL_NAND2X2 U9223 ( .A(n11030), .B(n10806), .Z(n10053) );
  HS65_LL_NAND2X2 U9224 ( .A(n10741), .B(n7989), .Z(n10941) );
  HS65_LL_NOR2X2 U9225 ( .A(n7969), .B(n10720), .Z(n10715) );
  HS65_LL_IVX2 U9226 ( .A(n10715), .Z(n10807) );
  HS65_LL_NAND2X2 U9227 ( .A(n10956), .B(n7989), .Z(n11057) );
  HS65_LL_NAND3X2 U9228 ( .A(n10941), .B(n10807), .C(n11057), .Z(n13369) );
  HS65_LL_NAND2X2 U9229 ( .A(n7958), .B(n7967), .Z(n10742) );
  HS65_LL_NAND2X2 U9230 ( .A(n10742), .B(n7955), .Z(n13375) );
  HS65_LL_NOR2X2 U9231 ( .A(n10060), .B(n7959), .Z(n10620) );
  HS65_LL_IVX2 U9232 ( .A(n10060), .Z(n10740) );
  HS65_LL_NAND2X2 U9233 ( .A(n10740), .B(n7956), .Z(n13367) );
  HS65_LL_NAND2X2 U9234 ( .A(n11022), .B(n13367), .Z(n10722) );
  HS65_LL_NOR2X2 U9235 ( .A(n10620), .B(n10722), .Z(n10746) );
  HS65_LL_NAND4ABX3 U9236 ( .A(n13369), .B(n13375), .C(n10746), .D(n10739), 
        .Z(n7957) );
  HS65_LL_NOR3X1 U9237 ( .A(n10624), .B(n10053), .C(n7957), .Z(n11046) );
  HS65_LL_NOR2X2 U9238 ( .A(n10056), .B(n7959), .Z(n13383) );
  HS65_LL_IVX2 U9239 ( .A(n10637), .Z(n11033) );
  HS65_LL_NOR2X2 U9240 ( .A(n13383), .B(n11033), .Z(n10618) );
  HS65_LL_NOR2X2 U9241 ( .A(n10824), .B(n10629), .Z(n10736) );
  HS65_LL_NAND2X2 U9242 ( .A(n7958), .B(n10956), .Z(n10626) );
  HS65_LL_IVX2 U9243 ( .A(n10626), .Z(n10619) );
  HS65_LL_NOR2X2 U9244 ( .A(n10736), .B(n10619), .Z(n7960) );
  HS65_LL_NOR2X2 U9245 ( .A(n11025), .B(n7983), .Z(n10825) );
  HS65_LL_NOR2X2 U9246 ( .A(n10060), .B(n11025), .Z(n13366) );
  HS65_LL_NOR2X2 U9247 ( .A(n7959), .B(n7983), .Z(n10833) );
  HS65_LL_NOR2X2 U9248 ( .A(n13366), .B(n10833), .Z(n11035) );
  HS65_LL_OAI21X2 U9249 ( .A(sa12[7]), .B(n13391), .C(n11035), .Z(n13382) );
  HS65_LL_NOR4ABX2 U9250 ( .A(n7960), .B(n10614), .C(n10825), .D(n13382), .Z(
        n7962) );
  HS65_LL_NOR2X2 U9251 ( .A(n7969), .B(n10824), .Z(n10061) );
  HS65_LL_NOR2X2 U9252 ( .A(n11024), .B(n10629), .Z(n10639) );
  HS65_LL_NOR2X2 U9253 ( .A(n11025), .B(n10960), .Z(n11050) );
  HS65_LL_NOR2X2 U9254 ( .A(n7979), .B(n11050), .Z(n10069) );
  HS65_LL_NAND2X2 U9255 ( .A(n7985), .B(n10612), .Z(n7981) );
  HS65_LL_NAND4ABX3 U9256 ( .A(n10061), .B(n10639), .C(n10069), .D(n7981), .Z(
        n10814) );
  HS65_LL_IVX2 U9257 ( .A(n10052), .Z(n7966) );
  HS65_LL_NOR2X2 U9258 ( .A(n10060), .B(n7966), .Z(n11043) );
  HS65_LL_NAND2AX4 U9259 ( .A(n11043), .B(n10948), .Z(n7961) );
  HS65_LL_NOR4ABX2 U9260 ( .A(n10618), .B(n7962), .C(n10814), .D(n7961), .Z(
        n7996) );
  HS65_LL_NAND2X2 U9261 ( .A(sa12[4]), .B(sa12[2]), .Z(n10756) );
  HS65_LL_NOR2X2 U9262 ( .A(sa12[1]), .B(n10735), .Z(n11048) );
  HS65_LL_NAND3X2 U9263 ( .A(sa12[6]), .B(n10641), .C(n7963), .Z(n10815) );
  HS65_LL_IVX2 U9264 ( .A(n10815), .Z(n10609) );
  HS65_LL_IVX2 U9265 ( .A(n10941), .Z(n10934) );
  HS65_LL_NOR2AX3 U9266 ( .A(n11022), .B(n10825), .Z(n7965) );
  HS65_LL_NOR2X2 U9267 ( .A(n7969), .B(n7983), .Z(n10743) );
  HS65_LL_NOR2X2 U9268 ( .A(n10743), .B(n10930), .Z(n10731) );
  HS65_LL_NOR2X2 U9269 ( .A(n10056), .B(n10629), .Z(n13365) );
  HS65_LL_IVX2 U9270 ( .A(n13365), .Z(n7964) );
  HS65_LL_NAND2X2 U9271 ( .A(n10740), .B(n10641), .Z(n10826) );
  HS65_LL_NAND2X2 U9272 ( .A(n7964), .B(n10826), .Z(n10054) );
  HS65_LL_NOR2AX3 U9273 ( .A(n10731), .B(n10054), .Z(n11055) );
  HS65_LL_NAND4ABX3 U9274 ( .A(n13400), .B(n10934), .C(n7965), .D(n11055), .Z(
        n7978) );
  HS65_LL_NOR2X2 U9275 ( .A(n7966), .B(n7968), .Z(n11060) );
  HS65_LL_NAND2X2 U9276 ( .A(n7967), .B(n7989), .Z(n10617) );
  HS65_LL_NOR2X2 U9277 ( .A(n7969), .B(n7968), .Z(n10607) );
  HS65_LL_NOR4ABX2 U9278 ( .A(n10948), .B(n10617), .C(n10620), .D(n10607), .Z(
        n7971) );
  HS65_LL_NAND2X2 U9279 ( .A(n10641), .B(n7970), .Z(n11045) );
  HS65_LL_NAND3AX3 U9280 ( .A(n11060), .B(n7971), .C(n11045), .Z(n13379) );
  HS65_LL_NOR2X2 U9281 ( .A(n7972), .B(n10824), .Z(n10954) );
  HS65_LL_NAND3X2 U9282 ( .A(sa12[5]), .B(sa12[3]), .C(n7973), .Z(n10613) );
  HS65_LL_NAND2X2 U9283 ( .A(n7975), .B(n7974), .Z(n10831) );
  HS65_LL_NAND3AX3 U9284 ( .A(n10954), .B(n10613), .C(n10831), .Z(n7976) );
  HS65_LL_NOR3X1 U9285 ( .A(n13379), .B(n10608), .C(n7976), .Z(n10713) );
  HS65_LL_NAND4ABX3 U9286 ( .A(n10609), .B(n7978), .C(n10713), .D(n7977), .Z(
        n10966) );
  HS65_LL_NAND2X2 U9287 ( .A(n10614), .B(n10807), .Z(n10634) );
  HS65_LL_NOR2X2 U9288 ( .A(n7979), .B(n10634), .Z(n10644) );
  HS65_LL_NAND4ABX3 U9289 ( .A(n11064), .B(n10966), .C(n10644), .D(n13367), 
        .Z(n7994) );
  HS65_LL_NOR2X2 U9290 ( .A(sa12[4]), .B(sa12[2]), .Z(n13401) );
  HS65_LL_IVX2 U9291 ( .A(n10607), .Z(n7980) );
  HS65_LL_NAND2X2 U9292 ( .A(n10609), .B(n10623), .Z(n13384) );
  HS65_LL_NOR4ABX2 U9293 ( .A(n7980), .B(n13384), .C(n10811), .D(n10931), .Z(
        n13371) );
  HS65_LL_NOR2X2 U9294 ( .A(n10060), .B(n10051), .Z(n10734) );
  HS65_LL_NOR4ABX2 U9295 ( .A(n11057), .B(n7981), .C(n11043), .D(n10734), .Z(
        n7982) );
  HS65_LL_NOR4ABX2 U9296 ( .A(n13371), .B(n7982), .C(n10073), .D(n13377), .Z(
        n10823) );
  HS65_LL_NOR3X1 U9297 ( .A(n7985), .B(n7984), .C(n7983), .Z(n7986) );
  HS65_LL_NOR3X1 U9298 ( .A(n13366), .B(n13365), .C(n7986), .Z(n10943) );
  HS65_LL_IVX2 U9299 ( .A(n10061), .Z(n11037) );
  HS65_LL_IVX2 U9300 ( .A(n10831), .Z(n7987) );
  HS65_LL_NAND2X2 U9301 ( .A(sa12[5]), .B(n7987), .Z(n11042) );
  HS65_LL_OAI21X2 U9302 ( .A(n10720), .B(n7988), .C(n11042), .Z(n10936) );
  HS65_LL_AOI12X2 U9303 ( .A(n7989), .B(n10641), .C(n11060), .Z(n10726) );
  HS65_LL_NAND3X2 U9304 ( .A(n10726), .B(n7990), .C(n10637), .Z(n10837) );
  HS65_LL_NOR4ABX2 U9305 ( .A(n10943), .B(n11037), .C(n10936), .D(n10837), .Z(
        n7992) );
  HS65_LL_NOR2X2 U9306 ( .A(sa12[2]), .B(n7991), .Z(n11068) );
  HS65_LL_IVX2 U9307 ( .A(n11068), .Z(n13407) );
  HS65_LL_AOI13X2 U9308 ( .A(n10065), .B(n10823), .C(n7992), .D(n13407), .Z(
        n7993) );
  HS65_LL_CBI4I6X2 U9309 ( .A(n11048), .B(n7994), .C(n13401), .D(n7993), .Z(
        n7995) );
  HS65_LL_CBI4I1X3 U9310 ( .A(n11046), .B(n7996), .C(n10756), .D(n7995), .Z(
        n7997) );
  HS65_LL_CBI4I6X2 U9311 ( .A(n7999), .B(n7998), .C(n13410), .D(n7997), .Z(
        n15266) );
  HS65_LL_MUXI21X2 U9312 ( .D0(n15360), .D1(w1[14]), .S0(n15266), .Z(n8000) );
  HS65_LLS_XOR3X2 U9313 ( .A(n12148), .B(n14957), .C(n8000), .Z(n8001) );
  HS65_LL_MUXI21X2 U9314 ( .D0(n15361), .D1(n14983), .S0(n8001), .Z(n8002) );
  HS65_LL_IVX2 U9315 ( .A(ld_r), .Z(n11557) );
  HS65_LL_BFX4 U9316 ( .A(n11557), .Z(n14808) );
  HS65_LL_MUX31X4 U9317 ( .D0(w1[14]), .D1(n15360), .D2(n8002), .S0(
        text_in_r[78]), .S1(n14808), .Z(N184) );
  HS65_LL_BFX4 U9318 ( .A(n15806), .Z(n15843) );
  HS65_LL_IVX2 U9319 ( .A(w3[29]), .Z(n15242) );
  HS65_LL_IVX2 U9320 ( .A(w2[29]), .Z(n15571) );
  HS65_LL_IVX2 U9321 ( .A(w1[29]), .Z(n15128) );
  HS65_LL_IVX2 U9322 ( .A(w0[29]), .Z(n15526) );
  HS65_LL_NAND2X2 U9323 ( .A(n10383), .B(n8003), .Z(n10334) );
  HS65_LL_NOR4ABX2 U9324 ( .A(n8004), .B(n8024), .C(n8038), .D(n10495), .Z(
        n10380) );
  HS65_LL_NAND4ABX3 U9325 ( .A(n10468), .B(n10334), .C(n10380), .D(n10494), 
        .Z(n8017) );
  HS65_LL_NOR2X2 U9326 ( .A(n8006), .B(n8005), .Z(n8010) );
  HS65_LL_IVX2 U9327 ( .A(n10506), .Z(n8007) );
  HS65_LL_OAI21X2 U9328 ( .A(n10523), .B(n8018), .C(n8007), .Z(n10391) );
  HS65_LL_NOR2X2 U9329 ( .A(n10456), .B(n10492), .Z(n10317) );
  HS65_LL_NAND3X2 U9330 ( .A(n10317), .B(n10522), .C(n8019), .Z(n8008) );
  HS65_LL_NOR3X1 U9331 ( .A(n10493), .B(n10316), .C(n8008), .Z(n10462) );
  HS65_LL_NAND2X2 U9332 ( .A(n8012), .B(n8023), .Z(n10405) );
  HS65_LL_NAND3X2 U9333 ( .A(n10462), .B(n8029), .C(n10405), .Z(n8009) );
  HS65_LL_NOR3X1 U9334 ( .A(n8010), .B(n10391), .C(n8009), .Z(n15074) );
  HS65_LL_NOR2X2 U9335 ( .A(n15077), .B(n10321), .Z(n10392) );
  HS65_LL_NAND4ABX3 U9336 ( .A(n10376), .B(n8011), .C(n15074), .D(n10392), .Z(
        n8016) );
  HS65_LL_AOI12X2 U9337 ( .A(n8012), .B(n8026), .C(n10511), .Z(n10386) );
  HS65_LL_NAND2AX4 U9338 ( .A(n10374), .B(n8013), .Z(n15066) );
  HS65_LL_NOR4ABX2 U9339 ( .A(n10386), .B(n8014), .C(n10365), .D(n15066), .Z(
        n10437) );
  HS65_LL_NOR3X1 U9340 ( .A(n8015), .B(n10340), .C(n10490), .Z(n10526) );
  HS65_LL_NAND4ABX3 U9341 ( .A(n8017), .B(n8016), .C(n10437), .D(n10526), .Z(
        n8052) );
  HS65_LL_NOR2X2 U9342 ( .A(n15048), .B(n8018), .Z(n10370) );
  HS65_LL_NAND2X2 U9343 ( .A(n10367), .B(n8019), .Z(n10390) );
  HS65_LL_NOR3X1 U9344 ( .A(n10370), .B(n10312), .C(n10390), .Z(n10454) );
  HS65_LL_NOR2X2 U9345 ( .A(w3[17]), .B(w3[22]), .Z(n10423) );
  HS65_LL_NOR2X2 U9346 ( .A(n15691), .B(n8020), .Z(n10500) );
  HS65_LL_NOR2X2 U9347 ( .A(n10419), .B(n10500), .Z(n10418) );
  HS65_LL_NOR2X2 U9348 ( .A(n10406), .B(n8033), .Z(n10425) );
  HS65_LL_NAND3AX3 U9349 ( .A(n8021), .B(n10418), .C(n10425), .Z(n10473) );
  HS65_LL_CBI4I6X2 U9350 ( .A(n10423), .B(n8023), .C(n8022), .D(n10473), .Z(
        n8025) );
  HS65_LL_NOR4ABX2 U9351 ( .A(n8025), .B(n8024), .C(n15062), .D(n10321), .Z(
        n10319) );
  HS65_LL_AOI12X2 U9352 ( .A(n8026), .B(n10422), .C(n10365), .Z(n10323) );
  HS65_LL_NAND2X2 U9353 ( .A(n10323), .B(n8027), .Z(n10313) );
  HS65_LL_NOR4ABX2 U9354 ( .A(n10319), .B(n8028), .C(n10443), .D(n10313), .Z(
        n8030) );
  HS65_LL_NAND2X2 U9355 ( .A(n8029), .B(n10486), .Z(n10336) );
  HS65_LL_NOR4ABX2 U9356 ( .A(n8030), .B(n10517), .C(n10468), .D(n10336), .Z(
        n8031) );
  HS65_LL_NAND3X2 U9357 ( .A(n10363), .B(n10454), .C(n8031), .Z(n8051) );
  HS65_LL_NOR4ABX2 U9358 ( .A(n8034), .B(n10446), .C(n8033), .D(n8032), .Z(
        n10333) );
  HS65_LL_NOR2X2 U9359 ( .A(n8036), .B(n8035), .Z(n10410) );
  HS65_LL_NOR2X2 U9360 ( .A(n10485), .B(n10484), .Z(n8037) );
  HS65_LL_NAND4ABX3 U9361 ( .A(n8038), .B(n10464), .C(n8037), .D(n10361), .Z(
        n8039) );
  HS65_LL_NOR4ABX2 U9362 ( .A(n8040), .B(n8046), .C(n10410), .D(n8039), .Z(
        n8041) );
  HS65_LL_NAND3X2 U9363 ( .A(n10333), .B(n8042), .C(n8041), .Z(n8050) );
  HS65_LL_NOR2X2 U9364 ( .A(n10364), .B(n10320), .Z(n10338) );
  HS65_LL_NAND2X2 U9365 ( .A(n10338), .B(n10315), .Z(n10521) );
  HS65_LL_NOR3AX2 U9366 ( .A(n10494), .B(n10410), .C(n10312), .Z(n10346) );
  HS65_LL_IVX2 U9367 ( .A(n10500), .Z(n10384) );
  HS65_LL_NOR4ABX2 U9368 ( .A(n10384), .B(n10516), .C(n10484), .D(n15068), .Z(
        n8044) );
  HS65_LL_NOR2X2 U9369 ( .A(n15046), .B(n8043), .Z(n10382) );
  HS65_LL_NOR4ABX2 U9370 ( .A(n8045), .B(n8044), .C(n10343), .D(n10382), .Z(
        n10537) );
  HS65_LL_NOR4ABX2 U9371 ( .A(n10537), .B(n8046), .C(n10365), .D(n10391), .Z(
        n8047) );
  HS65_LL_NAND4ABX3 U9372 ( .A(n10521), .B(n8048), .C(n10346), .D(n8047), .Z(
        n8049) );
  HS65_LL_IVX2 U9373 ( .A(n10535), .Z(n15082) );
  HS65_LL_MX41X4 U9374 ( .D0(n8052), .S0(n15088), .D1(n8051), .S1(n15086), 
        .D2(n8050), .S2(n15084), .D3(n8049), .S3(n15082), .Z(n8053) );
  HS65_LLS_XOR3X2 U9375 ( .A(\u0/rcon [29]), .B(n15526), .C(n8053), .Z(n10359)
         );
  HS65_LL_MUXI21X2 U9376 ( .D0(n15128), .D1(w1[29]), .S0(n10359), .Z(n10483)
         );
  HS65_LL_MUXI21X2 U9377 ( .D0(n15571), .D1(w2[29]), .S0(n10483), .Z(n11618)
         );
  HS65_LL_MUX31X4 U9378 ( .D0(n15242), .D1(w3[29]), .D2(key[29]), .S0(n11618), 
        .S1(n15783), .Z(\u0/N269 ) );
  HS65_LL_IVX2 U9379 ( .A(w2[19]), .Z(n15332) );
  HS65_LL_IVX2 U9380 ( .A(sa20[1]), .Z(n8784) );
  HS65_LL_NOR3X1 U9381 ( .A(sa20[7]), .B(sa20[6]), .C(n8784), .Z(n8058) );
  HS65_LL_IVX2 U9382 ( .A(n8058), .Z(n8083) );
  HS65_LL_IVX2 U9383 ( .A(sa20[5]), .Z(n8078) );
  HS65_LL_NAND3X2 U9384 ( .A(sa20[3]), .B(sa20[0]), .C(n8078), .Z(n8076) );
  HS65_LL_NOR2X2 U9385 ( .A(n8083), .B(n8076), .Z(n8800) );
  HS65_LL_IVX2 U9386 ( .A(sa20[7]), .Z(n8088) );
  HS65_LL_NOR3X1 U9387 ( .A(sa20[1]), .B(sa20[6]), .C(n8088), .Z(n8070) );
  HS65_LL_IVX2 U9388 ( .A(n8070), .Z(n8059) );
  HS65_LL_NOR2X2 U9389 ( .A(n8059), .B(n8076), .Z(n12340) );
  HS65_LL_IVX2 U9390 ( .A(sa20[6]), .Z(n8057) );
  HS65_LL_NOR2X2 U9391 ( .A(n8057), .B(sa20[7]), .Z(n8322) );
  HS65_LL_NAND2X2 U9392 ( .A(n8784), .B(n8322), .Z(n8242) );
  HS65_LL_NAND3X2 U9393 ( .A(sa20[5]), .B(sa20[3]), .C(sa20[0]), .Z(n8237) );
  HS65_LL_NOR2X2 U9394 ( .A(n8242), .B(n8237), .Z(n8776) );
  HS65_LL_NOR2X2 U9395 ( .A(n12340), .B(n8776), .Z(n15386) );
  HS65_LL_NAND2AX4 U9396 ( .A(n8800), .B(n15386), .Z(n8239) );
  HS65_LL_NOR3X1 U9397 ( .A(sa20[1]), .B(sa20[7]), .C(sa20[6]), .Z(n9036) );
  HS65_LL_IVX2 U9398 ( .A(n9036), .Z(n8067) );
  HS65_LL_NOR2X2 U9399 ( .A(n8067), .B(n8076), .Z(n12341) );
  HS65_LL_NAND3X2 U9400 ( .A(sa20[1]), .B(sa20[7]), .C(sa20[6]), .Z(n8085) );
  HS65_LL_IVX2 U9401 ( .A(n8085), .Z(n8054) );
  HS65_LL_NOR2X2 U9402 ( .A(sa20[3]), .B(sa20[0]), .Z(n8055) );
  HS65_LL_NAND2X2 U9403 ( .A(n8055), .B(n8078), .Z(n8091) );
  HS65_LL_IVX2 U9404 ( .A(n8091), .Z(n8318) );
  HS65_LL_NAND2X2 U9405 ( .A(n8054), .B(n8318), .Z(n12303) );
  HS65_LL_IVX2 U9406 ( .A(n12303), .Z(n15380) );
  HS65_LL_NOR2X2 U9407 ( .A(n12341), .B(n15380), .Z(n8071) );
  HS65_LL_IVX2 U9408 ( .A(sa20[3]), .Z(n8077) );
  HS65_LL_NOR3AX2 U9409 ( .A(sa20[0]), .B(n8077), .C(n8059), .Z(n8774) );
  HS65_LL_NAND2X2 U9410 ( .A(n8774), .B(sa20[5]), .Z(n9035) );
  HS65_LL_NAND2X2 U9411 ( .A(n8071), .B(n9035), .Z(n15410) );
  HS65_LL_NAND2X2 U9412 ( .A(sa20[5]), .B(n8055), .Z(n8316) );
  HS65_LL_IVX2 U9413 ( .A(n8316), .Z(n8247) );
  HS65_LL_NAND2X2 U9414 ( .A(n8247), .B(n9036), .Z(n8794) );
  HS65_LL_IVX2 U9415 ( .A(n8794), .Z(n9055) );
  HS65_LL_AND2X4 U9416 ( .A(sa20[0]), .B(n8077), .Z(n8246) );
  HS65_LL_NAND2X2 U9417 ( .A(sa20[5]), .B(n8246), .Z(n8084) );
  HS65_LL_NOR2X2 U9418 ( .A(n8084), .B(n8085), .Z(n13040) );
  HS65_LL_NOR2X2 U9419 ( .A(n9055), .B(n13040), .Z(n9041) );
  HS65_LL_NOR2X2 U9420 ( .A(n8085), .B(n8237), .Z(n12301) );
  HS65_LL_NAND3X2 U9421 ( .A(sa20[7]), .B(sa20[6]), .C(n8784), .Z(n8092) );
  HS65_LL_NOR2X2 U9422 ( .A(n8092), .B(n8076), .Z(n15394) );
  HS65_LL_NOR2X2 U9423 ( .A(n12301), .B(n15394), .Z(n12332) );
  HS65_LL_NOR2X2 U9424 ( .A(n8084), .B(n8067), .Z(n8311) );
  HS65_LL_IVX2 U9425 ( .A(n8311), .Z(n12314) );
  HS65_LL_NAND3X2 U9426 ( .A(n9041), .B(n12332), .C(n12314), .Z(n8056) );
  HS65_LL_OR3X4 U9427 ( .A(n8239), .B(n15410), .C(n8056), .Z(n12299) );
  HS65_LL_NAND2X2 U9428 ( .A(n8078), .B(n8246), .Z(n8074) );
  HS65_LL_NAND3X2 U9429 ( .A(sa20[7]), .B(sa20[1]), .C(n8057), .Z(n8236) );
  HS65_LL_NOR2X2 U9430 ( .A(n8074), .B(n8236), .Z(n9044) );
  HS65_LL_IVX2 U9431 ( .A(n8084), .Z(n8073) );
  HS65_LL_NAND2X2 U9432 ( .A(sa20[1]), .B(n8322), .Z(n8317) );
  HS65_LL_IVX2 U9433 ( .A(n8317), .Z(n8066) );
  HS65_LL_NAND2X2 U9434 ( .A(n8073), .B(n8066), .Z(n8243) );
  HS65_LL_NOR2X2 U9435 ( .A(n8074), .B(n8085), .Z(n15384) );
  HS65_LL_NOR2X2 U9436 ( .A(n8316), .B(n8236), .Z(n12307) );
  HS65_LL_NOR2X2 U9437 ( .A(n15384), .B(n12307), .Z(n8080) );
  HS65_LL_NAND4ABX3 U9438 ( .A(n12299), .B(n9044), .C(n8243), .D(n8080), .Z(
        n8095) );
  HS65_LL_NOR2X2 U9439 ( .A(n8077), .B(sa20[0]), .Z(n9037) );
  HS65_LL_NAND2X2 U9440 ( .A(n9037), .B(n8078), .Z(n8344) );
  HS65_LL_NOR2X2 U9441 ( .A(n8059), .B(n8344), .Z(n13015) );
  HS65_LL_NAND2X2 U9442 ( .A(sa20[5]), .B(n9037), .Z(n8087) );
  HS65_LL_NOR2X2 U9443 ( .A(n8087), .B(n8067), .Z(n9065) );
  HS65_LL_OR2X4 U9444 ( .A(n13015), .B(n9065), .Z(n8773) );
  HS65_LL_NOR2X2 U9445 ( .A(n8087), .B(n8236), .Z(n8252) );
  HS65_LL_NOR2X2 U9446 ( .A(n8316), .B(n8092), .Z(n12324) );
  HS65_LL_NOR2X2 U9447 ( .A(n8252), .B(n12324), .Z(n8334) );
  HS65_LL_NOR2X2 U9448 ( .A(n8236), .B(n8076), .Z(n9075) );
  HS65_LL_NOR2X2 U9449 ( .A(n8344), .B(n8085), .Z(n9032) );
  HS65_LL_NOR2X2 U9450 ( .A(n9075), .B(n9032), .Z(n8064) );
  HS65_LL_IVX2 U9451 ( .A(n8236), .Z(n8330) );
  HS65_LL_NAND2X2 U9452 ( .A(n8318), .B(n8330), .Z(n8782) );
  HS65_LL_NOR2X2 U9453 ( .A(n8059), .B(n8316), .Z(n12315) );
  HS65_LL_IVX2 U9454 ( .A(n8074), .Z(n8062) );
  HS65_LL_NAND2X2 U9455 ( .A(n8058), .B(n8062), .Z(n8244) );
  HS65_LL_NOR2X2 U9456 ( .A(n8074), .B(n8092), .Z(n8313) );
  HS65_LL_IVX2 U9457 ( .A(n8313), .Z(n13017) );
  HS65_LL_AND2X4 U9458 ( .A(n8244), .B(n13017), .Z(n15381) );
  HS65_LL_NOR2X2 U9459 ( .A(n8317), .B(n8344), .Z(n8235) );
  HS65_LL_NOR2X2 U9460 ( .A(n8059), .B(n8087), .Z(n13034) );
  HS65_LL_NOR2X2 U9461 ( .A(n8235), .B(n13034), .Z(n8771) );
  HS65_LL_NOR2X2 U9462 ( .A(n8087), .B(n8242), .Z(n9074) );
  HS65_LL_NOR2X2 U9463 ( .A(n8074), .B(n8317), .Z(n8331) );
  HS65_LL_NOR2X2 U9464 ( .A(n9074), .B(n8331), .Z(n9058) );
  HS65_LL_NOR2X2 U9465 ( .A(n8344), .B(n8067), .Z(n8329) );
  HS65_LL_IVX2 U9466 ( .A(n8329), .Z(n9072) );
  HS65_LL_NOR2X2 U9467 ( .A(n8084), .B(n8236), .Z(n12316) );
  HS65_LL_NOR2X2 U9468 ( .A(n8087), .B(n8085), .Z(n8786) );
  HS65_LL_NOR4ABX2 U9469 ( .A(n9058), .B(n9072), .C(n12316), .D(n8786), .Z(
        n8060) );
  HS65_LL_NAND3X2 U9470 ( .A(n15381), .B(n8771), .C(n8060), .Z(n15418) );
  HS65_LL_NOR4ABX2 U9471 ( .A(n8064), .B(n8782), .C(n12315), .D(n15418), .Z(
        n8061) );
  HS65_LL_NAND4ABX3 U9472 ( .A(n8095), .B(n8773), .C(n8334), .D(n8061), .Z(
        n8101) );
  HS65_LL_IVX2 U9473 ( .A(sa20[4]), .Z(n8097) );
  HS65_LL_NOR2X2 U9474 ( .A(sa20[2]), .B(n8097), .Z(n15416) );
  HS65_LL_NOR2X2 U9475 ( .A(n8084), .B(n8242), .Z(n8093) );
  HS65_LL_NOR2X2 U9476 ( .A(n9044), .B(n9055), .Z(n8230) );
  HS65_LL_NAND2X2 U9477 ( .A(n8070), .B(n8062), .Z(n12311) );
  HS65_LL_IVX2 U9478 ( .A(n8235), .Z(n9034) );
  HS65_LL_NAND2X2 U9479 ( .A(n8062), .B(n9036), .Z(n13032) );
  HS65_LL_NAND2X2 U9480 ( .A(n9034), .B(n13032), .Z(n8338) );
  HS65_LL_NOR4ABX2 U9481 ( .A(n8230), .B(n12311), .C(n8773), .D(n8338), .Z(
        n8063) );
  HS65_LL_NAND4ABX3 U9482 ( .A(n8093), .B(n8786), .C(n8064), .D(n8063), .Z(
        n8336) );
  HS65_LL_NOR2X2 U9483 ( .A(n8344), .B(n8236), .Z(n12323) );
  HS65_LL_NOR2X2 U9484 ( .A(n8085), .B(n8076), .Z(n8339) );
  HS65_LL_NOR2X2 U9485 ( .A(n12323), .B(n8339), .Z(n8328) );
  HS65_LL_NOR2X2 U9486 ( .A(n8317), .B(n8237), .Z(n13014) );
  HS65_LL_NOR2X2 U9487 ( .A(n8252), .B(n13014), .Z(n15397) );
  HS65_LL_NAND2X2 U9488 ( .A(n8070), .B(n8318), .Z(n8319) );
  HS65_LL_IVX2 U9489 ( .A(n15384), .Z(n8314) );
  HS65_LL_NOR2X2 U9490 ( .A(n8083), .B(n8344), .Z(n15407) );
  HS65_LL_NOR4ABX2 U9491 ( .A(n8319), .B(n8314), .C(n12340), .D(n15407), .Z(
        n8065) );
  HS65_LL_AND3X4 U9492 ( .A(n8328), .B(n15397), .C(n8065), .Z(n15374) );
  HS65_LL_NOR2X2 U9493 ( .A(n8092), .B(n8237), .Z(n12308) );
  HS65_LL_NAND2X2 U9494 ( .A(n8066), .B(n8318), .Z(n15382) );
  HS65_LL_IVX2 U9495 ( .A(n15382), .Z(n8248) );
  HS65_LL_NOR2X2 U9496 ( .A(n12308), .B(n8248), .Z(n9059) );
  HS65_LL_NOR2X2 U9497 ( .A(n8067), .B(n8237), .Z(n8778) );
  HS65_LL_NOR2X2 U9498 ( .A(n8778), .B(n9074), .Z(n12297) );
  HS65_LL_NOR2X2 U9499 ( .A(n8083), .B(n8091), .Z(n8787) );
  HS65_LL_IVX2 U9500 ( .A(n8787), .Z(n13035) );
  HS65_LL_NOR3X1 U9501 ( .A(sa20[7]), .B(sa20[6]), .C(n8084), .Z(n8781) );
  HS65_LL_NOR4ABX2 U9502 ( .A(n12297), .B(n13035), .C(n15380), .D(n8781), .Z(
        n8068) );
  HS65_LL_NOR2X2 U9503 ( .A(n8083), .B(n8087), .Z(n8249) );
  HS65_LL_NOR4ABX2 U9504 ( .A(n9059), .B(n8068), .C(n15394), .D(n8249), .Z(
        n8069) );
  HS65_LL_NAND3AX3 U9505 ( .A(n8336), .B(n15374), .C(n8069), .Z(n8100) );
  HS65_LL_NOR2X2 U9506 ( .A(sa20[2]), .B(sa20[4]), .Z(n13020) );
  HS65_LL_NAND2X2 U9507 ( .A(sa20[6]), .B(n8784), .Z(n8089) );
  HS65_LL_NAND2X2 U9508 ( .A(n8073), .B(n8070), .Z(n8793) );
  HS65_LL_OAI112X1 U9509 ( .A(n8237), .B(n8089), .C(n8793), .D(n9072), .Z(
        n8082) );
  HS65_LL_NOR3AX2 U9510 ( .A(n8071), .B(n8252), .C(n8339), .Z(n9049) );
  HS65_LL_NOR2X2 U9511 ( .A(n8242), .B(n8076), .Z(n12306) );
  HS65_LL_NOR2X2 U9512 ( .A(n8093), .B(n12315), .Z(n8775) );
  HS65_LL_IVX2 U9513 ( .A(n8092), .Z(n8072) );
  HS65_LL_NAND2X2 U9514 ( .A(n8073), .B(n8072), .Z(n9068) );
  HS65_LL_IVX2 U9515 ( .A(n9068), .Z(n8255) );
  HS65_LL_NOR2AX3 U9516 ( .A(n8775), .B(n8255), .Z(n15373) );
  HS65_LL_NOR2X2 U9517 ( .A(n12340), .B(n12301), .Z(n9062) );
  HS65_LL_NOR2X2 U9518 ( .A(n8074), .B(n8242), .Z(n15395) );
  HS65_LL_IVX2 U9519 ( .A(n8344), .Z(n8785) );
  HS65_LL_NAND3X2 U9520 ( .A(sa20[7]), .B(sa20[6]), .C(n8785), .Z(n12302) );
  HS65_LL_NOR2X2 U9521 ( .A(sa20[1]), .B(n12302), .Z(n8251) );
  HS65_LL_NOR2X2 U9522 ( .A(n15395), .B(n8251), .Z(n8796) );
  HS65_LL_NAND3X2 U9523 ( .A(n15373), .B(n9062), .C(n8796), .Z(n8075) );
  HS65_LL_NOR3X1 U9524 ( .A(n8778), .B(n12324), .C(n8075), .Z(n13047) );
  HS65_LL_NOR2X2 U9525 ( .A(n13015), .B(n8311), .Z(n8250) );
  HS65_LL_IVX2 U9526 ( .A(n8243), .Z(n8779) );
  HS65_LL_NOR3X1 U9527 ( .A(sa20[7]), .B(n8784), .C(n8076), .Z(n12300) );
  HS65_LL_NAND2X2 U9528 ( .A(sa20[6]), .B(n12300), .Z(n9050) );
  HS65_LL_NOR3X1 U9529 ( .A(n8078), .B(n8077), .C(n8083), .Z(n9067) );
  HS65_LL_NAND2X2 U9530 ( .A(sa20[0]), .B(n9067), .Z(n13023) );
  HS65_LL_NOR3X1 U9531 ( .A(sa20[3]), .B(sa20[0]), .C(n8083), .Z(n12310) );
  HS65_LL_NAND2X2 U9532 ( .A(sa20[5]), .B(n12310), .Z(n15392) );
  HS65_LL_NAND3X2 U9533 ( .A(n9050), .B(n13023), .C(n15392), .Z(n15376) );
  HS65_LL_NOR3X1 U9534 ( .A(n8779), .B(n13034), .C(n15376), .Z(n8079) );
  HS65_LL_NAND3X2 U9535 ( .A(n13047), .B(n8250), .C(n8079), .Z(n8234) );
  HS65_LL_NOR4ABX2 U9536 ( .A(n8080), .B(n13035), .C(n12306), .D(n8234), .Z(
        n8081) );
  HS65_LL_NAND4ABX3 U9537 ( .A(n9032), .B(n8082), .C(n9049), .D(n8081), .Z(
        n8099) );
  HS65_LL_AND2X4 U9538 ( .A(sa20[2]), .B(sa20[4]), .Z(n15408) );
  HS65_LL_NOR2X2 U9539 ( .A(n8084), .B(n8083), .Z(n9061) );
  HS65_LL_IVX2 U9540 ( .A(n9061), .Z(n8343) );
  HS65_LL_NAND2X2 U9541 ( .A(n8343), .B(n12311), .Z(n8257) );
  HS65_LL_NOR2X2 U9542 ( .A(n8317), .B(n8087), .Z(n9071) );
  HS65_LL_IVX2 U9543 ( .A(n9071), .Z(n9045) );
  HS65_LL_NAND2X2 U9544 ( .A(n9045), .B(n8793), .Z(n9060) );
  HS65_LL_IVX2 U9545 ( .A(n15395), .Z(n13036) );
  HS65_LL_NOR2X2 U9546 ( .A(n8316), .B(n8085), .Z(n8324) );
  HS65_LL_NOR2X2 U9547 ( .A(n8324), .B(n8329), .Z(n8340) );
  HS65_LL_NAND4ABX3 U9548 ( .A(n8235), .B(n12308), .C(n13036), .D(n8340), .Z(
        n8086) );
  HS65_LL_NOR3X1 U9549 ( .A(n8257), .B(n9060), .C(n8086), .Z(n8241) );
  HS65_LL_NAND2X2 U9550 ( .A(n8319), .B(n8244), .Z(n12330) );
  HS65_LL_NOR3X1 U9551 ( .A(sa20[6]), .B(n8784), .C(n8091), .Z(n9038) );
  HS65_LL_NOR2X2 U9552 ( .A(n8088), .B(n8087), .Z(n8259) );
  HS65_LL_NOR2AX3 U9553 ( .A(n8259), .B(n8089), .Z(n8312) );
  HS65_LL_OR3X4 U9554 ( .A(n8312), .B(n13015), .C(n8252), .Z(n8090) );
  HS65_LL_NOR3X1 U9555 ( .A(n12330), .B(n9038), .C(n8090), .Z(n13027) );
  HS65_LL_NOR2X2 U9556 ( .A(n8092), .B(n8091), .Z(n9073) );
  HS65_LL_IVX2 U9557 ( .A(n8093), .Z(n8315) );
  HS65_LL_NAND4ABX3 U9558 ( .A(n12316), .B(n9073), .C(n8315), .D(n13017), .Z(
        n8094) );
  HS65_LL_NOR3X1 U9559 ( .A(n8095), .B(n15376), .C(n8094), .Z(n8096) );
  HS65_LL_NAND3X2 U9560 ( .A(n8241), .B(n13027), .C(n8096), .Z(n8098) );
  HS65_LL_NAND2X2 U9561 ( .A(n8097), .B(sa20[2]), .Z(n13045) );
  HS65_LL_IVX2 U9562 ( .A(n13045), .Z(n15400) );
  HS65_LL_MX41X4 U9563 ( .D0(n8101), .S0(n15416), .D1(n8100), .S1(n13020), 
        .D2(n8099), .S2(n15408), .D3(n8098), .S3(n15400), .Z(n15423) );
  HS65_LL_IVX2 U9564 ( .A(n15423), .Z(n15424) );
  HS65_LL_NOR2X2 U9565 ( .A(sa13[7]), .B(sa13[6]), .Z(n9000) );
  HS65_LL_IVX2 U9566 ( .A(sa13[1]), .Z(n8808) );
  HS65_LL_NAND2X2 U9567 ( .A(n9000), .B(n8808), .Z(n8816) );
  HS65_LL_NOR2X2 U9568 ( .A(sa13[0]), .B(sa13[3]), .Z(n8989) );
  HS65_LL_NAND2X2 U9569 ( .A(sa13[5]), .B(n8989), .Z(n8814) );
  HS65_LL_NOR2X2 U9570 ( .A(n8816), .B(n8814), .Z(n8287) );
  HS65_LL_NAND3X2 U9571 ( .A(sa13[7]), .B(sa13[6]), .C(sa13[1]), .Z(n8114) );
  HS65_LL_IVX2 U9572 ( .A(sa13[3]), .Z(n8296) );
  HS65_LL_AND2X4 U9573 ( .A(sa13[0]), .B(n8296), .Z(n8818) );
  HS65_LL_NAND2X2 U9574 ( .A(sa13[5]), .B(n8818), .Z(n8832) );
  HS65_LL_NOR2X2 U9575 ( .A(n8114), .B(n8832), .Z(n14515) );
  HS65_LL_NOR2X2 U9576 ( .A(n8287), .B(n14515), .Z(n9015) );
  HS65_LL_NAND2X2 U9577 ( .A(sa13[0]), .B(sa13[3]), .Z(n8990) );
  HS65_LL_NOR2X2 U9578 ( .A(sa13[5]), .B(n8990), .Z(n8281) );
  HS65_LL_NOR2X2 U9579 ( .A(n8816), .B(n8832), .Z(n8840) );
  HS65_LL_AOI12X2 U9580 ( .A(n9000), .B(n8281), .C(n8840), .Z(n8104) );
  HS65_LL_IVX2 U9581 ( .A(n8990), .Z(n8664) );
  HS65_LL_NAND2X2 U9582 ( .A(sa13[5]), .B(n8664), .Z(n14521) );
  HS65_LL_IVX2 U9583 ( .A(sa13[6]), .Z(n15282) );
  HS65_LL_NOR2X2 U9584 ( .A(n15282), .B(sa13[7]), .Z(n8105) );
  HS65_LL_NAND2X2 U9585 ( .A(n8105), .B(n8808), .Z(n8279) );
  HS65_LL_NOR2X2 U9586 ( .A(n14521), .B(n8279), .Z(n8641) );
  HS65_LL_IVX2 U9587 ( .A(n8281), .Z(n15281) );
  HS65_LL_NAND3X2 U9588 ( .A(sa13[6]), .B(sa13[7]), .C(n8808), .Z(n8111) );
  HS65_LL_NOR2X2 U9589 ( .A(n15281), .B(n8111), .Z(n12278) );
  HS65_LL_NOR2X2 U9590 ( .A(n8641), .B(n12278), .Z(n8102) );
  HS65_LL_NAND3X2 U9591 ( .A(sa13[7]), .B(n15282), .C(n8808), .Z(n8831) );
  HS65_LL_NOR2X2 U9592 ( .A(n14521), .B(n8831), .Z(n15289) );
  HS65_LL_IVX2 U9593 ( .A(n15289), .Z(n9007) );
  HS65_LL_IVX2 U9594 ( .A(sa13[5]), .Z(n8996) );
  HS65_LL_NAND2X2 U9595 ( .A(n8989), .B(n8996), .Z(n8266) );
  HS65_LL_NOR2X2 U9596 ( .A(n8114), .B(n8266), .Z(n15317) );
  HS65_LL_IVX2 U9597 ( .A(n8114), .Z(n8663) );
  HS65_LL_IVX2 U9598 ( .A(n14521), .Z(n8298) );
  HS65_LL_NAND2X2 U9599 ( .A(n8663), .B(n8298), .Z(n8810) );
  HS65_LL_IVX2 U9600 ( .A(n8831), .Z(n8817) );
  HS65_LL_NAND2X2 U9601 ( .A(n8281), .B(n8817), .Z(n15304) );
  HS65_LL_NAND2X2 U9602 ( .A(n8810), .B(n15304), .Z(n8998) );
  HS65_LL_NOR4ABX2 U9603 ( .A(n8102), .B(n9007), .C(n15317), .D(n8998), .Z(
        n8103) );
  HS65_LL_NAND3X2 U9604 ( .A(n9015), .B(n8104), .C(n8103), .Z(n12265) );
  HS65_LL_NAND2X2 U9605 ( .A(n8996), .B(n8818), .Z(n8267) );
  HS65_LL_IVX2 U9606 ( .A(n8267), .Z(n8118) );
  HS65_LL_AND2X4 U9607 ( .A(sa13[7]), .B(n15282), .Z(n8116) );
  HS65_LL_NAND2X2 U9608 ( .A(sa13[1]), .B(n8116), .Z(n8988) );
  HS65_LL_IVX2 U9609 ( .A(n8988), .Z(n8297) );
  HS65_LL_NAND2X2 U9610 ( .A(n8118), .B(n8297), .Z(n9025) );
  HS65_LL_IVX2 U9611 ( .A(n8832), .Z(n8108) );
  HS65_LL_NAND3X2 U9612 ( .A(sa13[1]), .B(n8105), .C(n8108), .Z(n15296) );
  HS65_LL_NAND2X2 U9613 ( .A(n9025), .B(n15296), .Z(n8299) );
  HS65_LL_NOR2X2 U9614 ( .A(n8814), .B(n8988), .Z(n8838) );
  HS65_LL_IVX2 U9615 ( .A(n8838), .Z(n12272) );
  HS65_LL_NOR2X2 U9616 ( .A(n8114), .B(n8267), .Z(n8653) );
  HS65_LL_IVX2 U9617 ( .A(n8653), .Z(n8645) );
  HS65_LL_NAND4ABX3 U9618 ( .A(n12265), .B(n8299), .C(n12272), .D(n8645), .Z(
        n8126) );
  HS65_LL_IVX2 U9619 ( .A(n8816), .Z(n8300) );
  HS65_LL_IVX2 U9620 ( .A(n8105), .Z(n14522) );
  HS65_LL_NOR2X2 U9621 ( .A(n8808), .B(n14522), .Z(n8286) );
  HS65_LL_NOR2X2 U9622 ( .A(sa13[0]), .B(n8296), .Z(n12264) );
  HS65_LL_NAND2X2 U9623 ( .A(n12264), .B(n8996), .Z(n9002) );
  HS65_LL_IVX2 U9624 ( .A(n9002), .Z(n8809) );
  HS65_LL_OAI21X2 U9625 ( .A(n8300), .B(n8286), .C(n8809), .Z(n8632) );
  HS65_LL_NAND2X2 U9626 ( .A(sa13[5]), .B(n12264), .Z(n8289) );
  HS65_LL_IVX2 U9627 ( .A(n8286), .Z(n8815) );
  HS65_LL_NOR2X2 U9628 ( .A(n8289), .B(n8815), .Z(n12247) );
  HS65_LL_NOR2X2 U9629 ( .A(n8831), .B(n8832), .Z(n15302) );
  HS65_LL_NOR2X2 U9630 ( .A(n12247), .B(n15302), .Z(n12250) );
  HS65_LL_NOR2X2 U9631 ( .A(n8114), .B(n8814), .Z(n8634) );
  HS65_LL_NOR3X1 U9632 ( .A(sa13[7]), .B(sa13[6]), .C(n8808), .Z(n12263) );
  HS65_LL_NAND2X2 U9633 ( .A(n12263), .B(n8108), .Z(n8273) );
  HS65_LL_NAND2X2 U9634 ( .A(n8118), .B(n8817), .Z(n12280) );
  HS65_LL_NAND2X2 U9635 ( .A(n8273), .B(n12280), .Z(n8270) );
  HS65_LL_IVX2 U9636 ( .A(n8279), .Z(n8630) );
  HS65_LL_NAND2X2 U9637 ( .A(n8630), .B(n8118), .Z(n15278) );
  HS65_LL_IVX2 U9638 ( .A(n8111), .Z(n8112) );
  HS65_LL_NAND2X2 U9639 ( .A(n8298), .B(n8112), .Z(n8822) );
  HS65_LL_NAND2X2 U9640 ( .A(n15278), .B(n8822), .Z(n9022) );
  HS65_LL_NOR3X1 U9641 ( .A(n8634), .B(n8270), .C(n9022), .Z(n8106) );
  HS65_LL_NAND3X2 U9642 ( .A(n8632), .B(n12250), .C(n8106), .Z(n8302) );
  HS65_LL_NOR2X2 U9643 ( .A(n8289), .B(n8111), .Z(n8280) );
  HS65_LL_IVX2 U9644 ( .A(n12263), .Z(n8995) );
  HS65_LL_NOR2X2 U9645 ( .A(n8995), .B(n8267), .Z(n12240) );
  HS65_LL_NOR2X2 U9646 ( .A(n8280), .B(n12240), .Z(n15298) );
  HS65_LL_NAND2X2 U9647 ( .A(n8809), .B(n8817), .Z(n14520) );
  HS65_LL_IVX2 U9648 ( .A(n8266), .Z(n8629) );
  HS65_LL_NAND2X2 U9649 ( .A(n8629), .B(n8817), .Z(n12239) );
  HS65_LL_NAND2X2 U9650 ( .A(n8629), .B(n12263), .Z(n8805) );
  HS65_LL_NAND2X2 U9651 ( .A(n12239), .B(n8805), .Z(n8107) );
  HS65_LL_NAND2X2 U9652 ( .A(n8629), .B(n8297), .Z(n8842) );
  HS65_LL_IVX2 U9653 ( .A(n8289), .Z(n8117) );
  HS65_LL_NAND2X2 U9654 ( .A(n8117), .B(n8297), .Z(n15305) );
  HS65_LL_NAND2X2 U9655 ( .A(n8842), .B(n15305), .Z(n8128) );
  HS65_LL_NOR4ABX2 U9656 ( .A(n15298), .B(n14520), .C(n8107), .D(n8128), .Z(
        n14530) );
  HS65_LL_NAND2X2 U9657 ( .A(n8630), .B(n8108), .Z(n8659) );
  HS65_LL_NAND2X2 U9658 ( .A(n8629), .B(n8112), .Z(n8992) );
  HS65_LL_NOR2X2 U9659 ( .A(n8995), .B(n8814), .Z(n15280) );
  HS65_LL_NOR2X2 U9660 ( .A(n14521), .B(n8995), .Z(n14533) );
  HS65_LL_AOI112X2 U9661 ( .A(n8286), .B(n8281), .C(n15280), .D(n14533), .Z(
        n12269) );
  HS65_LL_IVX2 U9662 ( .A(n12269), .Z(n9014) );
  HS65_LL_NAND2X2 U9663 ( .A(n8118), .B(n8112), .Z(n15299) );
  HS65_LL_NOR2X2 U9664 ( .A(n8832), .B(n8988), .Z(n12248) );
  HS65_LL_IVX2 U9665 ( .A(n12248), .Z(n12279) );
  HS65_LL_NAND2X2 U9666 ( .A(n15299), .B(n12279), .Z(n8109) );
  HS65_LL_NOR4ABX2 U9667 ( .A(n8659), .B(n8992), .C(n9014), .D(n8109), .Z(
        n8110) );
  HS65_LL_NAND4ABX3 U9668 ( .A(n8126), .B(n8302), .C(n14530), .D(n8110), .Z(
        n8132) );
  HS65_LL_NOR2AX3 U9669 ( .A(sa13[2]), .B(sa13[4]), .Z(n15328) );
  HS65_LL_NOR2X2 U9670 ( .A(n15281), .B(n8279), .Z(n12258) );
  HS65_LL_IVX2 U9671 ( .A(n12258), .Z(n8295) );
  HS65_LL_NAND3X2 U9672 ( .A(n8295), .B(n12272), .C(n8822), .Z(n8654) );
  HS65_LL_NOR2X2 U9673 ( .A(n8114), .B(n9002), .Z(n12249) );
  HS65_LL_NAND3X2 U9674 ( .A(sa13[7]), .B(n8117), .C(n8808), .Z(n8269) );
  HS65_LL_NOR2X2 U9675 ( .A(sa13[6]), .B(n8269), .Z(n14514) );
  HS65_LL_IVX2 U9676 ( .A(n8814), .Z(n8285) );
  HS65_LL_NAND2X2 U9677 ( .A(n8285), .B(n8817), .Z(n8834) );
  HS65_LL_IVX2 U9678 ( .A(n8834), .Z(n12285) );
  HS65_LL_NOR2X2 U9679 ( .A(n8832), .B(n8111), .Z(n8987) );
  HS65_LL_NOR3AX2 U9680 ( .A(n8659), .B(n12285), .C(n8987), .Z(n8636) );
  HS65_LL_NAND2X2 U9681 ( .A(n12269), .B(n8636), .Z(n15321) );
  HS65_LL_NOR2AX3 U9682 ( .A(n14520), .B(n8840), .Z(n8277) );
  HS65_LL_NAND2X2 U9683 ( .A(n8285), .B(n8112), .Z(n12266) );
  HS65_LL_AND2X4 U9684 ( .A(n15278), .B(n12266), .Z(n8640) );
  HS65_LL_NAND2X2 U9685 ( .A(n8809), .B(n8112), .Z(n12276) );
  HS65_LL_NOR2X2 U9686 ( .A(n14521), .B(n8816), .Z(n12259) );
  HS65_LL_NOR4ABX2 U9687 ( .A(n8640), .B(n12276), .C(n12259), .D(n8998), .Z(
        n8635) );
  HS65_LL_NAND3X2 U9688 ( .A(n8277), .B(n8635), .C(n15296), .Z(n8113) );
  HS65_LL_NOR3X1 U9689 ( .A(n14514), .B(n15321), .C(n8113), .Z(n8293) );
  HS65_LL_NAND4ABX3 U9690 ( .A(n12249), .B(n8641), .C(n8645), .D(n8293), .Z(
        n8115) );
  HS65_LL_NAND2X2 U9691 ( .A(n8281), .B(n8300), .Z(n15291) );
  HS65_LL_OAI21X2 U9692 ( .A(n15281), .B(n8114), .C(n15305), .Z(n8122) );
  HS65_LL_NOR3AX2 U9693 ( .A(n15291), .B(n15317), .C(n8122), .Z(n9024) );
  HS65_LL_NAND2X2 U9694 ( .A(n8809), .B(n8300), .Z(n8993) );
  HS65_LL_IVX2 U9695 ( .A(n8993), .Z(n8643) );
  HS65_LL_IVX2 U9696 ( .A(n8805), .Z(n14516) );
  HS65_LL_NOR3X1 U9697 ( .A(n8643), .B(n14516), .C(n15302), .Z(n9012) );
  HS65_LL_NAND4ABX3 U9698 ( .A(n8654), .B(n8115), .C(n9024), .D(n9012), .Z(
        n8131) );
  HS65_LL_AND2X4 U9699 ( .A(sa13[2]), .B(sa13[4]), .Z(n15326) );
  HS65_LL_NAND2X2 U9700 ( .A(n8629), .B(n8286), .Z(n8652) );
  HS65_LL_NAND2X2 U9701 ( .A(n8652), .B(n8822), .Z(n9009) );
  HS65_LL_NOR2X2 U9702 ( .A(n9002), .B(n8815), .Z(n9006) );
  HS65_LL_NOR2X2 U9703 ( .A(n12249), .B(n9006), .Z(n8120) );
  HS65_LL_NAND2X2 U9704 ( .A(n8300), .B(n8117), .Z(n12237) );
  HS65_LL_NAND2X2 U9705 ( .A(n14520), .B(n12237), .Z(n8829) );
  HS65_LL_AOI112X2 U9706 ( .A(n8116), .B(n8118), .C(n8287), .D(n8829), .Z(
        n8119) );
  HS65_LL_NAND2X2 U9707 ( .A(n8663), .B(n8117), .Z(n15290) );
  HS65_LL_NAND2X2 U9708 ( .A(n15290), .B(n8659), .Z(n8282) );
  HS65_LL_NAND2X2 U9709 ( .A(n8300), .B(n8118), .Z(n9001) );
  HS65_LL_NAND2X2 U9710 ( .A(n8281), .B(n8297), .Z(n12260) );
  HS65_LL_NAND2X2 U9711 ( .A(n9001), .B(n12260), .Z(n14506) );
  HS65_LL_NOR4ABX2 U9712 ( .A(n8120), .B(n8119), .C(n8282), .D(n14506), .Z(
        n8649) );
  HS65_LL_NAND4ABX3 U9713 ( .A(n12259), .B(n9009), .C(n8273), .D(n8649), .Z(
        n8124) );
  HS65_LL_NOR2X2 U9714 ( .A(n14521), .B(n8815), .Z(n15279) );
  HS65_LL_NOR3X1 U9715 ( .A(sa13[6]), .B(n8808), .C(n9002), .Z(n8823) );
  HS65_LL_NOR2X2 U9716 ( .A(n15279), .B(n8823), .Z(n8639) );
  HS65_LL_NAND3X2 U9717 ( .A(n8639), .B(n12239), .C(n15304), .Z(n8121) );
  HS65_LL_NOR3X1 U9718 ( .A(n8653), .B(n8122), .C(n8121), .Z(n15318) );
  HS65_LL_NOR2X2 U9719 ( .A(n8995), .B(n8289), .Z(n8275) );
  HS65_LL_NOR2X2 U9720 ( .A(n8275), .B(n12278), .Z(n8291) );
  HS65_LL_NOR2X2 U9721 ( .A(n8279), .B(n8289), .Z(n12257) );
  HS65_LL_NOR4ABX2 U9722 ( .A(n8291), .B(n8805), .C(n12257), .D(n15317), .Z(
        n8123) );
  HS65_LL_NAND4ABX3 U9723 ( .A(n8840), .B(n8124), .C(n15318), .D(n8123), .Z(
        n8130) );
  HS65_LL_NOR2X2 U9724 ( .A(sa13[4]), .B(sa13[2]), .Z(n15324) );
  HS65_LL_NAND2X2 U9725 ( .A(n12266), .B(n12260), .Z(n8274) );
  HS65_LL_NOR4ABX2 U9726 ( .A(n8632), .B(n15290), .C(n12240), .D(n14514), .Z(
        n8125) );
  HS65_LL_NOR2X2 U9727 ( .A(n8267), .B(n8815), .Z(n8807) );
  HS65_LL_IVX2 U9728 ( .A(n8807), .Z(n12270) );
  HS65_LL_IVX2 U9729 ( .A(n12257), .Z(n14523) );
  HS65_LL_NAND2X2 U9730 ( .A(n12270), .B(n14523), .Z(n8997) );
  HS65_LL_NOR4ABX2 U9731 ( .A(n8125), .B(n15299), .C(n12248), .D(n8997), .Z(
        n15315) );
  HS65_LL_IVX2 U9732 ( .A(n12249), .Z(n9008) );
  HS65_LL_NOR4ABX2 U9733 ( .A(n9008), .B(n8834), .C(n8126), .D(n8829), .Z(
        n8127) );
  HS65_LL_NAND4ABX3 U9734 ( .A(n8274), .B(n8128), .C(n15315), .D(n8127), .Z(
        n8129) );
  HS65_LL_NOR2AX3 U9735 ( .A(sa13[4]), .B(sa13[2]), .Z(n15322) );
  HS65_LL_MX41X4 U9736 ( .D0(n8132), .S0(n15328), .D1(n8131), .S1(n15326), 
        .D2(n8130), .S2(n15324), .D3(n8129), .S3(n15322), .Z(n15607) );
  HS65_LL_MUXI21X2 U9737 ( .D0(n15424), .D1(n15423), .S0(n15607), .Z(n15630)
         );
  HS65_LL_IVX2 U9738 ( .A(sa31[7]), .Z(n8151) );
  HS65_LL_NOR2X2 U9739 ( .A(sa31[6]), .B(n8151), .Z(n8166) );
  HS65_LL_IVX2 U9740 ( .A(n8166), .Z(n8558) );
  HS65_LL_IVX2 U9741 ( .A(sa31[3]), .Z(n8138) );
  HS65_LL_IVX2 U9742 ( .A(sa31[0]), .Z(n8142) );
  HS65_LL_NOR2X2 U9743 ( .A(sa31[5]), .B(n8142), .Z(n8907) );
  HS65_LL_IVX2 U9744 ( .A(n8907), .Z(n8156) );
  HS65_LL_NOR2X2 U9745 ( .A(n8138), .B(n8156), .Z(n8740) );
  HS65_LL_IVX2 U9746 ( .A(sa31[1]), .Z(n12360) );
  HS65_LL_NAND2X2 U9747 ( .A(n8740), .B(n12360), .Z(n8903) );
  HS65_LL_NOR2X2 U9748 ( .A(n8558), .B(n8903), .Z(n12372) );
  HS65_LL_NAND2X2 U9749 ( .A(sa31[6]), .B(sa31[7]), .Z(n8733) );
  HS65_LL_NOR2X2 U9750 ( .A(n12360), .B(n8733), .Z(n8554) );
  HS65_LL_IVX2 U9751 ( .A(n8554), .Z(n8569) );
  HS65_LL_NAND3X2 U9752 ( .A(sa31[3]), .B(sa31[5]), .C(sa31[0]), .Z(n12375) );
  HS65_LL_NOR2X2 U9753 ( .A(n8569), .B(n12375), .Z(n13324) );
  HS65_LL_NOR2X2 U9754 ( .A(n12372), .B(n13324), .Z(n8557) );
  HS65_LL_NOR2X2 U9755 ( .A(n8733), .B(sa31[1]), .Z(n8147) );
  HS65_LL_NAND2X2 U9756 ( .A(sa31[5]), .B(n8142), .Z(n8585) );
  HS65_LL_NOR2X2 U9757 ( .A(sa31[3]), .B(n8585), .Z(n8563) );
  HS65_LL_NAND2X2 U9758 ( .A(n8147), .B(n8563), .Z(n8572) );
  HS65_LL_IVX2 U9759 ( .A(n8147), .Z(n8139) );
  HS65_LL_NOR2X2 U9760 ( .A(sa31[5]), .B(sa31[0]), .Z(n8910) );
  HS65_LL_NAND2X2 U9761 ( .A(sa31[3]), .B(n8910), .Z(n12369) );
  HS65_LL_NOR2X2 U9762 ( .A(n8139), .B(n12369), .Z(n12347) );
  HS65_LL_NAND3X2 U9763 ( .A(sa31[5]), .B(sa31[0]), .C(n8138), .Z(n8171) );
  HS65_LL_IVX2 U9764 ( .A(n8171), .Z(n8164) );
  HS65_LL_NAND3X2 U9765 ( .A(sa31[6]), .B(n12360), .C(n8151), .Z(n8738) );
  HS65_LL_IVX2 U9766 ( .A(n8738), .Z(n8134) );
  HS65_LL_NAND2X2 U9767 ( .A(n8164), .B(n8134), .Z(n8734) );
  HS65_LL_IVX2 U9768 ( .A(n8734), .Z(n8153) );
  HS65_LL_NOR2X2 U9769 ( .A(sa31[1]), .B(n8558), .Z(n8906) );
  HS65_LL_NAND2X2 U9770 ( .A(n8906), .B(n8563), .Z(n13076) );
  HS65_LL_NAND2X2 U9771 ( .A(n8147), .B(n8164), .Z(n13306) );
  HS65_LL_NAND2X2 U9772 ( .A(n13076), .B(n13306), .Z(n8929) );
  HS65_LL_NOR2X2 U9773 ( .A(n8153), .B(n8929), .Z(n15456) );
  HS65_LL_NAND2X2 U9774 ( .A(n8907), .B(n8138), .Z(n8746) );
  HS65_LL_NOR2X2 U9775 ( .A(n8746), .B(n8738), .Z(n15472) );
  HS65_LL_IVX2 U9776 ( .A(n15472), .Z(n12348) );
  HS65_LL_IVX2 U9777 ( .A(sa31[6]), .Z(n12370) );
  HS65_LL_NAND3X2 U9778 ( .A(n12370), .B(n12360), .C(n8151), .Z(n8160) );
  HS65_LL_IVX2 U9779 ( .A(n8160), .Z(n8739) );
  HS65_LL_IVX2 U9780 ( .A(n12375), .Z(n8161) );
  HS65_LL_NAND2X2 U9781 ( .A(n8739), .B(n8161), .Z(n15483) );
  HS65_LL_NAND3X2 U9782 ( .A(n15456), .B(n12348), .C(n15483), .Z(n8133) );
  HS65_LL_NOR4ABX2 U9783 ( .A(n8557), .B(n8572), .C(n12347), .D(n8133), .Z(
        n13059) );
  HS65_LL_NAND2X2 U9784 ( .A(sa31[1]), .B(n8563), .Z(n8902) );
  HS65_LL_NOR2X2 U9785 ( .A(n8733), .B(n8902), .Z(n8753) );
  HS65_LL_NOR3X1 U9786 ( .A(sa31[3]), .B(sa31[5]), .C(sa31[0]), .Z(n8564) );
  HS65_LL_NAND2X2 U9787 ( .A(n8564), .B(n8906), .Z(n8749) );
  HS65_LL_NAND2X2 U9788 ( .A(n8134), .B(n8564), .Z(n13347) );
  HS65_LL_NAND2X2 U9789 ( .A(n8749), .B(n13347), .Z(n8913) );
  HS65_LL_NAND2X2 U9790 ( .A(n8739), .B(n8164), .Z(n12379) );
  HS65_LL_NAND3X2 U9791 ( .A(sa31[1]), .B(n12370), .C(n8151), .Z(n8143) );
  HS65_LL_IVX2 U9792 ( .A(n8564), .Z(n8169) );
  HS65_LL_NOR2X2 U9793 ( .A(n8143), .B(n8169), .Z(n8932) );
  HS65_LL_IVX2 U9794 ( .A(n8932), .Z(n8916) );
  HS65_LL_NAND2X2 U9795 ( .A(n12379), .B(n8916), .Z(n8586) );
  HS65_LL_NOR2X2 U9796 ( .A(n8160), .B(n12369), .Z(n8176) );
  HS65_LL_IVX2 U9797 ( .A(n8176), .Z(n13318) );
  HS65_LL_IVX2 U9798 ( .A(n8746), .Z(n8148) );
  HS65_LL_NAND2X2 U9799 ( .A(n8148), .B(n8739), .Z(n13060) );
  HS65_LL_NAND2X2 U9800 ( .A(n13318), .B(n13060), .Z(n13328) );
  HS65_LL_NAND3X2 U9801 ( .A(sa31[1]), .B(sa31[6]), .C(n8151), .Z(n8155) );
  HS65_LL_IVX2 U9802 ( .A(n8155), .Z(n8135) );
  HS65_LL_AND2X4 U9803 ( .A(n8740), .B(n8554), .Z(n8737) );
  HS65_LL_AOI12X2 U9804 ( .A(n8910), .B(n8135), .C(n8737), .Z(n8136) );
  HS65_LL_IVX2 U9805 ( .A(n8585), .Z(n8570) );
  HS65_LL_NAND2X2 U9806 ( .A(sa31[3]), .B(n8570), .Z(n8745) );
  HS65_LL_NOR3X1 U9807 ( .A(sa31[1]), .B(n8151), .C(n8745), .Z(n8728) );
  HS65_LL_NAND2X2 U9808 ( .A(sa31[6]), .B(n8728), .Z(n8565) );
  HS65_LL_NAND4ABX3 U9809 ( .A(n8586), .B(n13328), .C(n8136), .D(n8565), .Z(
        n8137) );
  HS65_LL_NOR3X1 U9810 ( .A(n8753), .B(n8913), .C(n8137), .Z(n12355) );
  HS65_LL_NAND2X2 U9811 ( .A(sa31[1]), .B(n8166), .Z(n12376) );
  HS65_LL_IVX2 U9812 ( .A(n12376), .Z(n8146) );
  HS65_LL_NAND2AX4 U9813 ( .A(n12369), .B(n8146), .Z(n13344) );
  HS65_LL_NOR2X2 U9814 ( .A(n8138), .B(n8143), .Z(n13303) );
  HS65_LL_NAND2X2 U9815 ( .A(n8910), .B(n13303), .Z(n15469) );
  HS65_LL_NAND2X2 U9816 ( .A(n13344), .B(n15469), .Z(n8582) );
  HS65_LL_NOR2X2 U9817 ( .A(n8738), .B(n12375), .Z(n13064) );
  HS65_LL_IVX2 U9818 ( .A(n13064), .Z(n8555) );
  HS65_LL_NOR2X2 U9819 ( .A(n8733), .B(n8903), .Z(n8940) );
  HS65_LL_IVX2 U9820 ( .A(n8940), .Z(n8899) );
  HS65_LL_NOR2X2 U9821 ( .A(n8139), .B(n8169), .Z(n13311) );
  HS65_LL_IVX2 U9822 ( .A(n13311), .Z(n8140) );
  HS65_LL_NAND3X2 U9823 ( .A(n8555), .B(n8899), .C(n8140), .Z(n15462) );
  HS65_LL_NOR2X2 U9824 ( .A(n8155), .B(n12375), .Z(n15471) );
  HS65_LL_NAND2X2 U9825 ( .A(sa31[5]), .B(sa31[0]), .Z(n8141) );
  HS65_LL_NOR3X1 U9826 ( .A(sa31[1]), .B(n12370), .C(n12369), .Z(n15458) );
  HS65_LL_NAND2X2 U9827 ( .A(n15458), .B(n8151), .Z(n8168) );
  HS65_LL_OAI21X2 U9828 ( .A(n12376), .B(n8141), .C(n8168), .Z(n8163) );
  HS65_LL_NAND3X2 U9829 ( .A(n8142), .B(sa31[3]), .C(n8554), .Z(n8159) );
  HS65_LL_IVX2 U9830 ( .A(n8143), .Z(n8909) );
  HS65_LL_NAND2X2 U9831 ( .A(n8164), .B(n8909), .Z(n12381) );
  HS65_LL_NOR2X2 U9832 ( .A(n8155), .B(n8745), .Z(n13310) );
  HS65_LL_NOR2AX3 U9833 ( .A(n12381), .B(n13310), .Z(n8560) );
  HS65_LL_NAND4ABX3 U9834 ( .A(n15471), .B(n8163), .C(n8159), .D(n8560), .Z(
        n8144) );
  HS65_LL_NOR3X1 U9835 ( .A(n8582), .B(n15462), .C(n8144), .Z(n8145) );
  HS65_LL_NAND3X2 U9836 ( .A(n13059), .B(n12355), .C(n8145), .Z(n8183) );
  HS65_LL_IVX2 U9837 ( .A(sa31[2]), .Z(n8179) );
  HS65_LL_NOR2X2 U9838 ( .A(sa31[4]), .B(n8179), .Z(n15478) );
  HS65_LL_NAND3X2 U9839 ( .A(sa31[1]), .B(n8740), .C(n8151), .Z(n12357) );
  HS65_LL_NOR2X2 U9840 ( .A(sa31[6]), .B(n12357), .Z(n12378) );
  HS65_LL_NOR2X2 U9841 ( .A(n8155), .B(n8169), .Z(n15484) );
  HS65_LL_IVX2 U9842 ( .A(n8906), .Z(n8170) );
  HS65_LL_NOR2X2 U9843 ( .A(n8746), .B(n8170), .Z(n8561) );
  HS65_LL_IVX2 U9844 ( .A(n8563), .Z(n12359) );
  HS65_LL_NOR2X2 U9845 ( .A(n8155), .B(n12359), .Z(n15493) );
  HS65_LL_NOR2X2 U9846 ( .A(n8561), .B(n15493), .Z(n12353) );
  HS65_LL_NOR2X2 U9847 ( .A(n8171), .B(n12376), .Z(n8934) );
  HS65_LL_IVX2 U9848 ( .A(n8934), .Z(n8741) );
  HS65_LL_NAND4ABX3 U9849 ( .A(n15484), .B(n8913), .C(n12353), .D(n8741), .Z(
        n13309) );
  HS65_LL_NOR2X2 U9850 ( .A(n8746), .B(n8569), .Z(n15485) );
  HS65_LL_IVX2 U9851 ( .A(n15485), .Z(n8724) );
  HS65_LL_NAND2X2 U9852 ( .A(n8148), .B(n8147), .Z(n8723) );
  HS65_LL_IVX2 U9853 ( .A(n8723), .Z(n13341) );
  HS65_LL_IVX2 U9854 ( .A(n12379), .Z(n8930) );
  HS65_LL_NAND2X2 U9855 ( .A(n8146), .B(n8740), .Z(n15482) );
  HS65_LL_NAND2X2 U9856 ( .A(n8147), .B(n8161), .Z(n12363) );
  HS65_LL_AND2X4 U9857 ( .A(n15482), .B(n12363), .Z(n13348) );
  HS65_LL_NOR2X2 U9858 ( .A(n8746), .B(n8155), .Z(n8933) );
  HS65_LL_NAND3X2 U9859 ( .A(sa31[6]), .B(n8740), .C(n12360), .Z(n15473) );
  HS65_LL_NOR2X2 U9860 ( .A(sa31[7]), .B(n15473), .Z(n8578) );
  HS65_LL_NAND2X2 U9861 ( .A(n8148), .B(n8909), .Z(n15486) );
  HS65_LL_IVX2 U9862 ( .A(n15486), .Z(n13346) );
  HS65_LL_NOR2X2 U9863 ( .A(n8155), .B(n8171), .Z(n8920) );
  HS65_LL_NOR2X2 U9864 ( .A(n13346), .B(n8920), .Z(n15470) );
  HS65_LL_IVX2 U9865 ( .A(n15471), .Z(n8583) );
  HS65_LL_NAND2X2 U9866 ( .A(n15470), .B(n8583), .Z(n8735) );
  HS65_LL_NAND4ABX3 U9867 ( .A(n15462), .B(n8735), .C(n13060), .D(n13306), .Z(
        n8149) );
  HS65_LL_NOR3X1 U9868 ( .A(n8933), .B(n8578), .C(n8149), .Z(n8150) );
  HS65_LL_OAI112X1 U9869 ( .A(n8151), .B(n8902), .C(n13348), .D(n8150), .Z(
        n13068) );
  HS65_LL_NAND4ABX3 U9870 ( .A(n8737), .B(n13068), .C(n8565), .D(n13344), .Z(
        n8152) );
  HS65_LL_NOR3X1 U9871 ( .A(n13341), .B(n8930), .C(n8152), .Z(n13321) );
  HS65_LL_NOR2X2 U9872 ( .A(n8746), .B(n12376), .Z(n13335) );
  HS65_LL_NOR2X2 U9873 ( .A(n8745), .B(n12376), .Z(n15489) );
  HS65_LL_NOR3X1 U9874 ( .A(n13335), .B(n15489), .C(n12347), .Z(n8742) );
  HS65_LL_NOR4ABX2 U9875 ( .A(n13321), .B(n8742), .C(n13324), .D(n8153), .Z(
        n8154) );
  HS65_LL_NAND4ABX3 U9876 ( .A(n12378), .B(n13309), .C(n8724), .D(n8154), .Z(
        n8182) );
  HS65_LL_NOR2X2 U9877 ( .A(sa31[4]), .B(sa31[2]), .Z(n15494) );
  HS65_LL_NOR2X2 U9878 ( .A(n8155), .B(n12369), .Z(n12362) );
  HS65_LL_NAND2X2 U9879 ( .A(n8570), .B(n8739), .Z(n8157) );
  HS65_LL_NOR2X2 U9880 ( .A(n12369), .B(n8170), .Z(n13066) );
  HS65_LL_IVX2 U9881 ( .A(n13066), .Z(n8571) );
  HS65_LL_NOR2X2 U9882 ( .A(n8156), .B(n12376), .Z(n13316) );
  HS65_LL_NAND2X2 U9883 ( .A(n8734), .B(n13060), .Z(n8919) );
  HS65_LL_NOR4ABX2 U9884 ( .A(n8157), .B(n8571), .C(n13316), .D(n8919), .Z(
        n8158) );
  HS65_LL_NAND4ABX3 U9885 ( .A(n12362), .B(n8561), .C(n8159), .D(n8158), .Z(
        n8590) );
  HS65_LL_NOR2X2 U9886 ( .A(n8160), .B(n8169), .Z(n13304) );
  HS65_LL_NOR2X2 U9887 ( .A(n8578), .B(n13304), .Z(n8911) );
  HS65_LL_NAND2X2 U9888 ( .A(n8911), .B(n8724), .Z(n13058) );
  HS65_LL_NOR2X2 U9889 ( .A(n12372), .B(n13311), .Z(n15487) );
  HS65_LL_NAND2X2 U9890 ( .A(n8161), .B(n8906), .Z(n12371) );
  HS65_LL_NOR4ABX2 U9891 ( .A(n12371), .B(n12381), .C(n8933), .D(n15493), .Z(
        n8162) );
  HS65_LL_NAND4ABX3 U9892 ( .A(n13058), .B(n8163), .C(n15487), .D(n8162), .Z(
        n13079) );
  HS65_LL_NAND2X2 U9893 ( .A(n8554), .B(n8164), .Z(n8931) );
  HS65_LL_NAND2X2 U9894 ( .A(n8931), .B(n12348), .Z(n13072) );
  HS65_LL_NOR4ABX2 U9895 ( .A(n8555), .B(n8572), .C(n15489), .D(n13072), .Z(
        n15463) );
  HS65_LL_IVX2 U9896 ( .A(n12357), .Z(n8172) );
  HS65_LL_NAND2X2 U9897 ( .A(sa31[6]), .B(n8172), .Z(n13336) );
  HS65_LL_NAND4ABX3 U9898 ( .A(n8176), .B(n8737), .C(n13336), .D(n13344), .Z(
        n8165) );
  HS65_LL_AOI12X2 U9899 ( .A(n8166), .B(n8563), .C(n8165), .Z(n8167) );
  HS65_LL_NAND4ABX3 U9900 ( .A(n8590), .B(n13079), .C(n15463), .D(n8167), .Z(
        n8181) );
  HS65_LL_NAND2X2 U9901 ( .A(sa31[4]), .B(sa31[2]), .Z(n15500) );
  HS65_LL_IVX2 U9902 ( .A(n15500), .Z(n13352) );
  HS65_LL_NAND2X2 U9903 ( .A(n8931), .B(n8168), .Z(n13322) );
  HS65_LL_NOR2X2 U9904 ( .A(n12376), .B(n8169), .Z(n12380) );
  HS65_LL_NOR2X2 U9905 ( .A(n12380), .B(n8737), .Z(n8173) );
  HS65_LL_NOR2X2 U9906 ( .A(n8171), .B(n8170), .Z(n12350) );
  HS65_LL_NOR3X1 U9907 ( .A(n8172), .B(n12350), .C(n13310), .Z(n8743) );
  HS65_LL_NAND3X2 U9908 ( .A(n8173), .B(n8743), .C(n12363), .Z(n8174) );
  HS65_LL_NOR2X2 U9909 ( .A(n13335), .B(n8920), .Z(n8559) );
  HS65_LL_AOI12X2 U9910 ( .A(n12369), .B(n12375), .C(n12376), .Z(n13315) );
  HS65_LL_NOR4ABX2 U9911 ( .A(n8559), .B(n8572), .C(n8932), .D(n13315), .Z(
        n8754) );
  HS65_LL_NAND4ABX3 U9912 ( .A(n8753), .B(n8174), .C(n8557), .D(n8754), .Z(
        n8178) );
  HS65_LL_NOR2X2 U9913 ( .A(n8569), .B(n8745), .Z(n8175) );
  HS65_LL_NOR3X1 U9914 ( .A(n8933), .B(n13341), .C(n8175), .Z(n8917) );
  HS65_LL_NOR2AX3 U9915 ( .A(n8728), .B(sa31[6]), .Z(n13305) );
  HS65_LL_NOR2X2 U9916 ( .A(n8176), .B(n12362), .Z(n8562) );
  HS65_LL_NOR2X2 U9917 ( .A(n8745), .B(n8738), .Z(n13067) );
  HS65_LL_IVX2 U9918 ( .A(n13067), .Z(n13337) );
  HS65_LL_NAND3X2 U9919 ( .A(n8562), .B(n8741), .C(n13337), .Z(n8177) );
  HS65_LL_NOR4ABX2 U9920 ( .A(n8917), .B(n15486), .C(n13305), .D(n8177), .Z(
        n15460) );
  HS65_LL_NAND4ABX3 U9921 ( .A(n13322), .B(n8178), .C(n15460), .D(n8911), .Z(
        n8180) );
  HS65_LL_NAND2X2 U9922 ( .A(sa31[4]), .B(n8179), .Z(n8574) );
  HS65_LL_IVX2 U9923 ( .A(n8574), .Z(n15503) );
  HS65_LL_MX41X4 U9924 ( .D0(n8183), .S0(n15478), .D1(n8182), .S1(n15494), 
        .D2(n8181), .S2(n13352), .D3(n8180), .S3(n15503), .Z(n14628) );
  HS65_LL_IVX2 U9925 ( .A(n14628), .Z(n15508) );
  HS65_LL_IVX2 U9926 ( .A(sa02[3]), .Z(n8674) );
  HS65_LL_NOR2X2 U9927 ( .A(sa02[0]), .B(n8674), .Z(n8612) );
  HS65_LL_IVX2 U9928 ( .A(sa02[5]), .Z(n8675) );
  HS65_LL_NAND2X2 U9929 ( .A(n8612), .B(n8675), .Z(n8203) );
  HS65_LL_IVX2 U9930 ( .A(sa02[6]), .Z(n8202) );
  HS65_LL_NOR2X2 U9931 ( .A(sa02[7]), .B(n8202), .Z(n8197) );
  HS65_LL_NAND2X2 U9932 ( .A(sa02[1]), .B(n8197), .Z(n8214) );
  HS65_LL_NOR2X2 U9933 ( .A(n8203), .B(n8214), .Z(n8973) );
  HS65_LL_NAND3X2 U9934 ( .A(sa02[7]), .B(sa02[1]), .C(n8202), .Z(n8952) );
  HS65_LL_IVX2 U9935 ( .A(sa02[0]), .Z(n8184) );
  HS65_LL_NOR2X2 U9936 ( .A(sa02[3]), .B(n8184), .Z(n8957) );
  HS65_LL_NAND2X2 U9937 ( .A(sa02[5]), .B(n8957), .Z(n8196) );
  HS65_LL_NOR2X2 U9938 ( .A(n8952), .B(n8196), .Z(n8696) );
  HS65_LL_NOR3X1 U9939 ( .A(sa02[1]), .B(sa02[7]), .C(sa02[6]), .Z(n8712) );
  HS65_LL_NAND2X2 U9940 ( .A(n8612), .B(n8712), .Z(n9129) );
  HS65_LL_NOR2X2 U9941 ( .A(sa02[5]), .B(n9129), .Z(n8691) );
  HS65_LL_IVX2 U9942 ( .A(n8612), .Z(n8185) );
  HS65_LL_NOR2X2 U9943 ( .A(n8675), .B(n8185), .Z(n8710) );
  HS65_LL_IVX2 U9944 ( .A(sa02[1]), .Z(n8875) );
  HS65_LL_NAND2X2 U9945 ( .A(n8197), .B(n8875), .Z(n8694) );
  HS65_LL_IVX2 U9946 ( .A(n8694), .Z(n8195) );
  HS65_LL_NAND2X2 U9947 ( .A(n8710), .B(n8195), .Z(n9123) );
  HS65_LL_NAND2X2 U9948 ( .A(n8957), .B(n8675), .Z(n8211) );
  HS65_LL_IVX2 U9949 ( .A(n8211), .Z(n8224) );
  HS65_LL_NAND3X2 U9950 ( .A(sa02[7]), .B(sa02[6]), .C(n8875), .Z(n8604) );
  HS65_LL_IVX2 U9951 ( .A(n8604), .Z(n8198) );
  HS65_LL_NAND2X2 U9952 ( .A(n8224), .B(n8198), .Z(n9083) );
  HS65_LL_NAND2X2 U9953 ( .A(n9123), .B(n9083), .Z(n14496) );
  HS65_LL_IVX2 U9954 ( .A(n8710), .Z(n8619) );
  HS65_LL_NAND3X2 U9955 ( .A(sa02[1]), .B(sa02[7]), .C(sa02[6]), .Z(n8599) );
  HS65_LL_NOR2X2 U9956 ( .A(n8619), .B(n8599), .Z(n15161) );
  HS65_LL_NOR2X2 U9957 ( .A(n8214), .B(n8211), .Z(n9124) );
  HS65_LL_NOR2X2 U9958 ( .A(n15161), .B(n9124), .Z(n8854) );
  HS65_LL_NOR2X2 U9959 ( .A(sa02[7]), .B(sa02[6]), .Z(n9112) );
  HS65_LL_NAND2X2 U9960 ( .A(sa02[1]), .B(n9112), .Z(n8673) );
  HS65_LL_NOR2X2 U9961 ( .A(n8673), .B(n8211), .Z(n9084) );
  HS65_LL_NAND2X2 U9962 ( .A(sa02[7]), .B(n8875), .Z(n8186) );
  HS65_LL_NOR2X2 U9963 ( .A(n8619), .B(n8186), .Z(n8192) );
  HS65_LL_IVX2 U9964 ( .A(n8192), .Z(n8692) );
  HS65_LL_NOR2X2 U9965 ( .A(sa02[6]), .B(n8692), .Z(n9099) );
  HS65_LL_NOR2X2 U9966 ( .A(n9084), .B(n9099), .Z(n8881) );
  HS65_LL_NAND4ABX3 U9967 ( .A(n8691), .B(n14496), .C(n8854), .D(n8881), .Z(
        n8187) );
  HS65_LL_NOR3X1 U9968 ( .A(n8973), .B(n8696), .C(n8187), .Z(n15147) );
  HS65_LL_NAND2X2 U9969 ( .A(sa02[0]), .B(sa02[3]), .Z(n8188) );
  HS65_LL_NOR2X2 U9970 ( .A(sa02[5]), .B(n8188), .Z(n8956) );
  HS65_LL_IVX2 U9971 ( .A(n8956), .Z(n8215) );
  HS65_LL_NAND3X2 U9972 ( .A(sa02[7]), .B(n8875), .C(n8202), .Z(n8209) );
  HS65_LL_NOR2X2 U9973 ( .A(n8215), .B(n8209), .Z(n9125) );
  HS65_LL_NAND3X2 U9974 ( .A(sa02[5]), .B(sa02[0]), .C(sa02[3]), .Z(n8953) );
  HS65_LL_NOR2X2 U9975 ( .A(n8599), .B(n8953), .Z(n9121) );
  HS65_LL_NOR2X2 U9976 ( .A(n9125), .B(n9121), .Z(n8602) );
  HS65_LL_NOR3X1 U9977 ( .A(sa02[7]), .B(n8875), .C(n8215), .Z(n8971) );
  HS65_LL_IVX2 U9978 ( .A(n8214), .Z(n8713) );
  HS65_LL_NAND2X2 U9979 ( .A(n8710), .B(n8713), .Z(n9082) );
  HS65_LL_IVX2 U9980 ( .A(n8209), .Z(n8958) );
  HS65_LL_NAND3X2 U9981 ( .A(sa02[5]), .B(n8958), .C(n8957), .Z(n15172) );
  HS65_LL_NAND2X2 U9982 ( .A(n9082), .B(n15172), .Z(n9118) );
  HS65_LL_NOR2X2 U9983 ( .A(n8971), .B(n9118), .Z(n8706) );
  HS65_LL_NOR2X2 U9984 ( .A(n8599), .B(n8215), .Z(n8698) );
  HS65_LL_NOR3X1 U9985 ( .A(sa02[0]), .B(sa02[3]), .C(n8675), .Z(n8711) );
  HS65_LL_IVX2 U9986 ( .A(n8711), .Z(n8695) );
  HS65_LL_NOR2X2 U9987 ( .A(n8599), .B(n8695), .Z(n8683) );
  HS65_LL_NOR4ABX2 U9988 ( .A(n8602), .B(n8706), .C(n8698), .D(n8683), .Z(
        n8190) );
  HS65_LL_NOR2X2 U9989 ( .A(n8599), .B(n8196), .Z(n8688) );
  HS65_LL_NOR3X1 U9990 ( .A(sa02[5]), .B(sa02[0]), .C(sa02[3]), .Z(n8598) );
  HS65_LL_IVX2 U9991 ( .A(n8598), .Z(n8621) );
  HS65_LL_NOR2X2 U9992 ( .A(n8952), .B(n8621), .Z(n8950) );
  HS65_LL_NOR2X2 U9993 ( .A(n8203), .B(n8694), .Z(n8945) );
  HS65_LL_NOR3X1 U9994 ( .A(n8688), .B(n8950), .C(n8945), .Z(n9133) );
  HS65_LL_NAND2X2 U9995 ( .A(n8956), .B(n8195), .Z(n15154) );
  HS65_LL_IVX2 U9996 ( .A(n15154), .Z(n8218) );
  HS65_LL_IVX2 U9997 ( .A(n8712), .Z(n8205) );
  HS65_LL_NOR2X2 U9998 ( .A(n8621), .B(n8205), .Z(n9098) );
  HS65_LL_NOR2X2 U9999 ( .A(n8218), .B(n9098), .Z(n14476) );
  HS65_LL_NOR2X2 U10000 ( .A(n8953), .B(n8604), .Z(n14475) );
  HS65_LL_NOR2X2 U10001 ( .A(n8214), .B(n8196), .Z(n8611) );
  HS65_LL_NOR2X2 U10002 ( .A(n8695), .B(n8604), .Z(n8871) );
  HS65_LL_NOR2X2 U10003 ( .A(n8952), .B(n8203), .Z(n8217) );
  HS65_LL_NOR2X2 U10004 ( .A(n8952), .B(n8211), .Z(n9092) );
  HS65_LL_NOR2X2 U10005 ( .A(n8952), .B(n8953), .Z(n8191) );
  HS65_LL_NOR3X1 U10006 ( .A(n8217), .B(n9092), .C(n8191), .Z(n9110) );
  HS65_LL_NOR2X2 U10007 ( .A(sa02[0]), .B(sa02[3]), .Z(n8223) );
  HS65_LL_IVX2 U10008 ( .A(n8673), .Z(n8709) );
  HS65_LL_NAND2X2 U10009 ( .A(n8223), .B(n8709), .Z(n8858) );
  HS65_LL_NOR2X2 U10010 ( .A(sa02[5]), .B(n8858), .Z(n14488) );
  HS65_LL_IVX2 U10011 ( .A(n14488), .Z(n8613) );
  HS65_LL_NAND4ABX3 U10012 ( .A(n8611), .B(n8871), .C(n9110), .D(n8613), .Z(
        n8678) );
  HS65_LL_NOR4ABX2 U10013 ( .A(n9133), .B(n14476), .C(n14475), .D(n8678), .Z(
        n8189) );
  HS65_LL_NAND3X2 U10014 ( .A(n15147), .B(n8190), .C(n8189), .Z(n8229) );
  HS65_LL_IVX2 U10015 ( .A(sa02[2]), .Z(n8201) );
  HS65_LL_NAND2X2 U10016 ( .A(n8201), .B(sa02[4]), .Z(n8891) );
  HS65_LL_IVX2 U10017 ( .A(n8891), .Z(n15186) );
  HS65_LL_NOR2X2 U10018 ( .A(n8215), .B(n8604), .Z(n15149) );
  HS65_LL_NOR2X2 U10019 ( .A(n8953), .B(n8694), .Z(n8851) );
  HS65_LL_NOR2X2 U10020 ( .A(n15149), .B(n8851), .Z(n8601) );
  HS65_LL_OAI21X2 U10021 ( .A(n8621), .B(n8604), .C(n8601), .Z(n15143) );
  HS65_LL_IVX2 U10022 ( .A(n8203), .Z(n9111) );
  HS65_LL_NAND3X2 U10023 ( .A(n8202), .B(sa02[1]), .C(n9111), .Z(n8975) );
  HS65_LL_IVX2 U10024 ( .A(n8975), .Z(n8617) );
  HS65_LL_NAND2X2 U10025 ( .A(sa02[1]), .B(sa02[6]), .Z(n8622) );
  HS65_LL_NOR2X2 U10026 ( .A(n8696), .B(n8191), .Z(n8210) );
  HS65_LL_NOR2X2 U10027 ( .A(n8673), .B(n8196), .Z(n8864) );
  HS65_LL_IVX2 U10028 ( .A(n8864), .Z(n9122) );
  HS65_LL_OAI112X1 U10029 ( .A(n8622), .B(n8619), .C(n8210), .D(n9122), .Z(
        n8194) );
  HS65_LL_NOR2X2 U10030 ( .A(n8953), .B(n8214), .Z(n8616) );
  HS65_LL_NOR2X2 U10031 ( .A(n8616), .B(n8945), .Z(n15150) );
  HS65_LL_NOR2X2 U10032 ( .A(n8973), .B(n8683), .Z(n8717) );
  HS65_LL_NAND2X2 U10033 ( .A(n8598), .B(n8195), .Z(n8868) );
  HS65_LL_NAND2X2 U10034 ( .A(n8598), .B(n8958), .Z(n8708) );
  HS65_LL_NAND2X2 U10035 ( .A(sa02[6]), .B(n8192), .Z(n8714) );
  HS65_LL_NAND2X2 U10036 ( .A(n8708), .B(n8714), .Z(n8596) );
  HS65_LL_NOR2X2 U10037 ( .A(n8621), .B(n8214), .Z(n9120) );
  HS65_LL_NOR2X2 U10038 ( .A(n8698), .B(n8691), .Z(n8213) );
  HS65_LL_NAND2X2 U10039 ( .A(n8957), .B(n8712), .Z(n8676) );
  HS65_LL_NAND4ABX3 U10040 ( .A(n14488), .B(n9120), .C(n8213), .D(n8676), .Z(
        n8193) );
  HS65_LL_NOR4ABX2 U10041 ( .A(n8717), .B(n8868), .C(n8596), .D(n8193), .Z(
        n8963) );
  HS65_LL_NAND4ABX3 U10042 ( .A(n8617), .B(n8194), .C(n15150), .D(n8963), .Z(
        n8200) );
  HS65_LL_NAND2X2 U10043 ( .A(n8224), .B(n8195), .Z(n9089) );
  HS65_LL_IVX2 U10044 ( .A(n9089), .Z(n15153) );
  HS65_LL_NOR2X2 U10045 ( .A(n8953), .B(n8205), .Z(n9100) );
  HS65_LL_NOR2X2 U10046 ( .A(n8203), .B(n8604), .Z(n8863) );
  HS65_LL_IVX2 U10047 ( .A(n8196), .Z(n8221) );
  HS65_LL_NAND2X2 U10048 ( .A(n8197), .B(n8221), .Z(n8853) );
  HS65_LL_NOR2X2 U10049 ( .A(sa02[1]), .B(n8853), .Z(n8605) );
  HS65_LL_NAND2X2 U10050 ( .A(n8958), .B(n8711), .Z(n8852) );
  HS65_LL_NAND2X2 U10051 ( .A(n8221), .B(n8198), .Z(n9101) );
  HS65_LL_NAND2X2 U10052 ( .A(n8852), .B(n9101), .Z(n8859) );
  HS65_LL_NOR2X2 U10053 ( .A(n8605), .B(n8859), .Z(n15141) );
  HS65_LL_NAND4ABX3 U10054 ( .A(n9100), .B(n8863), .C(n8602), .D(n15141), .Z(
        n8199) );
  HS65_LL_NOR3X1 U10055 ( .A(n8871), .B(n15153), .C(n8199), .Z(n14482) );
  HS65_LL_NOR2X2 U10056 ( .A(n8599), .B(n8203), .Z(n9088) );
  HS65_LL_IVX2 U10057 ( .A(n9088), .Z(n9116) );
  HS65_LL_NAND4ABX3 U10058 ( .A(n15143), .B(n8200), .C(n14482), .D(n9116), .Z(
        n8228) );
  HS65_LL_NOR2X2 U10059 ( .A(sa02[4]), .B(n8201), .Z(n15184) );
  HS65_LL_NOR2X2 U10060 ( .A(n8605), .B(n15161), .Z(n8701) );
  HS65_LL_NOR2X2 U10061 ( .A(n8205), .B(n8695), .Z(n9131) );
  HS65_LL_NOR2X2 U10062 ( .A(n8952), .B(n8215), .Z(n9097) );
  HS65_LL_NOR2X2 U10063 ( .A(n9131), .B(n9097), .Z(n15177) );
  HS65_LL_NOR2X2 U10064 ( .A(sa02[5]), .B(n8676), .Z(n14477) );
  HS65_LL_NAND2X2 U10065 ( .A(sa02[7]), .B(n8202), .Z(n8204) );
  HS65_LL_OAI22X1 U10066 ( .A(n8204), .B(n8211), .C(n8622), .D(n8203), .Z(
        n8206) );
  HS65_LL_NAND2X2 U10067 ( .A(n8958), .B(n9111), .Z(n8704) );
  HS65_LL_NOR2X2 U10068 ( .A(n8619), .B(n8205), .Z(n8855) );
  HS65_LL_IVX2 U10069 ( .A(n8855), .Z(n8883) );
  HS65_LL_NAND2X2 U10070 ( .A(n8704), .B(n8883), .Z(n8946) );
  HS65_LL_NOR3X1 U10071 ( .A(n14477), .B(n8206), .C(n8946), .Z(n8207) );
  HS65_LL_NAND3X2 U10072 ( .A(n8701), .B(n15177), .C(n8207), .Z(n8624) );
  HS65_LL_NOR2X2 U10073 ( .A(n8688), .B(n15153), .Z(n14490) );
  HS65_LL_IVX2 U10074 ( .A(n8851), .Z(n8208) );
  HS65_LL_NOR2X2 U10075 ( .A(n8952), .B(n8619), .Z(n15171) );
  HS65_LL_NOR4ABX2 U10076 ( .A(n14490), .B(n8208), .C(n15171), .D(n8871), .Z(
        n15163) );
  HS65_LL_NOR3AX2 U10077 ( .A(n14476), .B(n9125), .C(n9124), .Z(n8680) );
  HS65_LL_NOR2X2 U10078 ( .A(n8209), .B(n8953), .Z(n8877) );
  HS65_LL_NOR2X2 U10079 ( .A(n8864), .B(n8877), .Z(n8687) );
  HS65_LL_NOR2X2 U10080 ( .A(n8621), .B(n8604), .Z(n9106) );
  HS65_LL_NOR2X2 U10081 ( .A(n8214), .B(n8695), .Z(n8882) );
  HS65_LL_NOR4ABX2 U10082 ( .A(n8687), .B(n8210), .C(n9106), .D(n8882), .Z(
        n8212) );
  HS65_LL_NOR2X2 U10083 ( .A(n8599), .B(n8211), .Z(n14478) );
  HS65_LL_NOR4ABX2 U10084 ( .A(n8680), .B(n8212), .C(n14478), .D(n8945), .Z(
        n14466) );
  HS65_LL_NAND3X2 U10085 ( .A(n15163), .B(n8213), .C(n14466), .Z(n8216) );
  HS65_LL_NOR2X2 U10086 ( .A(n8952), .B(n8695), .Z(n8972) );
  HS65_LL_NOR2X2 U10087 ( .A(n8215), .B(n8214), .Z(n8686) );
  HS65_LL_NOR3X1 U10088 ( .A(n8217), .B(n8972), .C(n8686), .Z(n9093) );
  HS65_LL_NAND4ABX3 U10089 ( .A(n8624), .B(n8216), .C(n9093), .D(n8852), .Z(
        n8227) );
  HS65_LL_AND2X4 U10090 ( .A(sa02[4]), .B(sa02[2]), .Z(n15182) );
  HS65_LL_NOR2X2 U10091 ( .A(n9092), .B(n8863), .Z(n8702) );
  HS65_LL_IVX2 U10092 ( .A(n8702), .Z(n8961) );
  HS65_LL_NAND2X2 U10093 ( .A(n8956), .B(n8709), .Z(n8951) );
  HS65_LL_NOR2X2 U10094 ( .A(n9084), .B(n8611), .Z(n15165) );
  HS65_LL_IVX2 U10095 ( .A(n8616), .Z(n14493) );
  HS65_LL_NAND2X2 U10096 ( .A(n15165), .B(n14493), .Z(n14487) );
  HS65_LL_NOR2AX3 U10097 ( .A(n8714), .B(n14487), .Z(n8700) );
  HS65_LL_IVX2 U10098 ( .A(n8217), .Z(n8857) );
  HS65_LL_NOR3X1 U10099 ( .A(n9097), .B(n14475), .C(n8218), .Z(n8887) );
  HS65_LL_NOR4ABX2 U10100 ( .A(n8887), .B(n9101), .C(n14477), .D(n8683), .Z(
        n8220) );
  HS65_LL_IVX2 U10101 ( .A(n9124), .Z(n8219) );
  HS65_LL_NOR4ABX2 U10102 ( .A(n8220), .B(n8219), .C(n8972), .D(n15143), .Z(
        n14486) );
  HS65_LL_NAND2X2 U10103 ( .A(n8221), .B(n8712), .Z(n8862) );
  HS65_LL_NAND3X2 U10104 ( .A(n14486), .B(n8862), .C(n9083), .Z(n8222) );
  HS65_LL_NOR4ABX2 U10105 ( .A(n8700), .B(n8857), .C(n8698), .D(n8222), .Z(
        n9132) );
  HS65_LL_NAND4ABX3 U10106 ( .A(n15171), .B(n8961), .C(n8951), .D(n9132), .Z(
        n8225) );
  HS65_LL_NAND2X2 U10107 ( .A(n8223), .B(n8713), .Z(n15168) );
  HS65_LL_NAND2X2 U10108 ( .A(n8958), .B(n8224), .Z(n8684) );
  HS65_LL_NAND2X2 U10109 ( .A(n8684), .B(n8868), .Z(n8884) );
  HS65_LL_NOR4ABX2 U10110 ( .A(n8708), .B(n15168), .C(n8696), .D(n8884), .Z(
        n9102) );
  HS65_LL_NOR2X2 U10111 ( .A(n14478), .B(n9121), .Z(n8689) );
  HS65_LL_NAND4ABX3 U10112 ( .A(n8605), .B(n8225), .C(n9102), .D(n8689), .Z(
        n8226) );
  HS65_LL_NOR2X2 U10113 ( .A(sa02[2]), .B(sa02[4]), .Z(n15180) );
  HS65_LL_MX41X4 U10114 ( .D0(n8229), .S0(n15186), .D1(n8228), .S1(n15184), 
        .D2(n8227), .S2(n15182), .D3(n8226), .S3(n15180), .Z(n15189) );
  HS65_LL_MUXI21X2 U10115 ( .D0(n15508), .D1(n14628), .S0(n15189), .Z(n14847)
         );
  HS65_LL_AOI112X2 U10116 ( .A(n8247), .B(n8322), .C(n8252), .D(n8249), .Z(
        n8233) );
  HS65_LL_NOR3X1 U10117 ( .A(n8776), .B(n15394), .C(n9073), .Z(n15377) );
  HS65_LL_NAND4ABX3 U10118 ( .A(n8324), .B(n8312), .C(n8230), .D(n8319), .Z(
        n8231) );
  HS65_LL_NOR4ABX2 U10119 ( .A(n15377), .B(n9035), .C(n8786), .D(n8231), .Z(
        n8232) );
  HS65_LL_NAND4ABX3 U10120 ( .A(n8235), .B(n8234), .C(n8233), .D(n8232), .Z(
        n8265) );
  HS65_LL_NOR2X2 U10121 ( .A(n8237), .B(n8236), .Z(n8780) );
  HS65_LL_NOR3X1 U10122 ( .A(n9044), .B(n12323), .C(n8780), .Z(n9076) );
  HS65_LL_NOR4ABX2 U10123 ( .A(n9076), .B(n13035), .C(n8779), .D(n12324), .Z(
        n8326) );
  HS65_LL_NAND4ABX3 U10124 ( .A(n9067), .B(n15407), .C(n15373), .D(n8326), .Z(
        n8238) );
  HS65_LL_AOI12X2 U10125 ( .A(n8246), .B(n9036), .C(n8238), .Z(n15391) );
  HS65_LL_IVX2 U10126 ( .A(n12306), .Z(n15393) );
  HS65_LL_NAND2X2 U10127 ( .A(n9036), .B(n8318), .Z(n13016) );
  HS65_LL_NAND2X2 U10128 ( .A(n15393), .B(n13016), .Z(n13031) );
  HS65_LL_NOR4ABX2 U10129 ( .A(n9058), .B(n9049), .C(n8239), .D(n13031), .Z(
        n8240) );
  HS65_LL_NAND3X2 U10130 ( .A(n8241), .B(n15391), .C(n8240), .Z(n8264) );
  HS65_LL_NOR2X2 U10131 ( .A(n12300), .B(n9060), .Z(n13038) );
  HS65_LL_IVX2 U10132 ( .A(n8242), .Z(n13019) );
  HS65_LL_NAND2X2 U10133 ( .A(n8244), .B(n8243), .Z(n8258) );
  HS65_LL_AOI12X2 U10134 ( .A(sa20[6]), .B(n8259), .C(n8258), .Z(n15405) );
  HS65_LL_NOR2AX3 U10135 ( .A(n8782), .B(n8339), .Z(n8323) );
  HS65_LL_NAND3AX3 U10136 ( .A(n13014), .B(n15405), .C(n8323), .Z(n8245) );
  HS65_LL_AOI12X2 U10137 ( .A(n8246), .B(n13019), .C(n8245), .Z(n12318) );
  HS65_LL_NAND2X2 U10138 ( .A(n13038), .B(n12318), .Z(n8772) );
  HS65_LL_NAND2X2 U10139 ( .A(n13019), .B(n8247), .Z(n12317) );
  HS65_LL_IVX2 U10140 ( .A(n12317), .Z(n9033) );
  HS65_LL_NOR2X2 U10141 ( .A(n12341), .B(n9033), .Z(n8795) );
  HS65_LL_NOR2X2 U10142 ( .A(n12316), .B(n8248), .Z(n12322) );
  HS65_LL_AOI12X2 U10143 ( .A(n9037), .B(n9036), .C(n9061), .Z(n12305) );
  HS65_LL_NAND3X2 U10144 ( .A(n8795), .B(n12322), .C(n12305), .Z(n13028) );
  HS65_LL_NOR3X1 U10145 ( .A(n9075), .B(n8249), .C(n12324), .Z(n12296) );
  HS65_LL_NAND2X2 U10146 ( .A(n12303), .B(n13016), .Z(n13039) );
  HS65_LL_NOR4ABX2 U10147 ( .A(n8250), .B(n12296), .C(n8776), .D(n13039), .Z(
        n9057) );
  HS65_LL_NOR3X1 U10148 ( .A(n8252), .B(n9044), .C(n8251), .Z(n8320) );
  HS65_LL_NOR4ABX2 U10149 ( .A(n8320), .B(n9068), .C(n15394), .D(n12315), .Z(
        n8253) );
  HS65_LL_NAND4ABX3 U10150 ( .A(n8772), .B(n13028), .C(n9057), .D(n8253), .Z(
        n8263) );
  HS65_LL_NOR2X2 U10151 ( .A(n15407), .B(n13031), .Z(n12294) );
  HS65_LL_NOR2X2 U10152 ( .A(n9071), .B(n9032), .Z(n13025) );
  HS65_LL_NAND2X2 U10153 ( .A(n8314), .B(n15392), .Z(n13029) );
  HS65_LL_NOR3X1 U10154 ( .A(n12301), .B(n8313), .C(n13029), .Z(n8254) );
  HS65_LL_NAND3X2 U10155 ( .A(n12294), .B(n13025), .C(n8254), .Z(n8798) );
  HS65_LL_IVX2 U10156 ( .A(n15394), .Z(n12325) );
  HS65_LL_IVX2 U10157 ( .A(n8331), .Z(n8788) );
  HS65_LL_NAND2X2 U10158 ( .A(n12325), .B(n8788), .Z(n12309) );
  HS65_LL_OR2X4 U10159 ( .A(n8324), .B(n8255), .Z(n12321) );
  HS65_LL_IVX2 U10160 ( .A(n8778), .Z(n9066) );
  HS65_LL_NAND3X2 U10161 ( .A(n9035), .B(n9050), .C(n9066), .Z(n8256) );
  HS65_LL_NOR3X1 U10162 ( .A(n8257), .B(n12321), .C(n8256), .Z(n8792) );
  HS65_LL_NOR2X2 U10163 ( .A(n13014), .B(n8258), .Z(n8308) );
  HS65_LL_NAND4ABX3 U10164 ( .A(n13040), .B(n12309), .C(n8792), .D(n8308), .Z(
        n8261) );
  HS65_LL_NOR3X1 U10165 ( .A(sa20[7]), .B(sa20[6]), .C(n8344), .Z(n9053) );
  HS65_LL_OAI21X2 U10166 ( .A(n8259), .B(n9053), .C(n8784), .Z(n8260) );
  HS65_LL_NAND4ABX3 U10167 ( .A(n8798), .B(n8261), .C(n9049), .D(n8260), .Z(
        n8262) );
  HS65_LL_MX41X4 U10168 ( .D0(n8265), .S0(n13020), .D1(n8264), .S1(n15416), 
        .D2(n8263), .S2(n15408), .D3(n8262), .S3(n15400), .Z(n15649) );
  HS65_LL_IVX2 U10169 ( .A(n15649), .Z(n15648) );
  HS65_LL_NAND2X2 U10170 ( .A(sa13[7]), .B(sa13[6]), .Z(n8288) );
  HS65_LL_IVX2 U10171 ( .A(n8810), .Z(n8658) );
  HS65_LL_NOR3X1 U10172 ( .A(n12249), .B(n8658), .C(n12258), .Z(n12277) );
  HS65_LL_NOR2X2 U10173 ( .A(n8266), .B(n8816), .Z(n14526) );
  HS65_LL_NOR2X2 U10174 ( .A(n9002), .B(n8995), .Z(n15293) );
  HS65_LL_NOR2X2 U10175 ( .A(n14526), .B(n15293), .Z(n14512) );
  HS65_LL_OAI112X1 U10176 ( .A(n8288), .B(n8267), .C(n12277), .D(n14512), .Z(
        n8268) );
  HS65_LL_NOR3X1 U10177 ( .A(n12247), .B(n15280), .C(n8268), .Z(n8828) );
  HS65_LL_NOR2X2 U10178 ( .A(n15279), .B(n12240), .Z(n15300) );
  HS65_LL_NAND2X2 U10179 ( .A(n15300), .B(n15296), .Z(n8655) );
  HS65_LL_NOR4ABX2 U10180 ( .A(n12270), .B(n8269), .C(n12278), .D(n8655), .Z(
        n8272) );
  HS65_LL_NOR2X2 U10181 ( .A(n8634), .B(n8987), .Z(n12271) );
  HS65_LL_AOI12X2 U10182 ( .A(n8286), .B(n8281), .C(n12259), .Z(n9020) );
  HS65_LL_NAND4ABX3 U10183 ( .A(n15289), .B(n8270), .C(n12271), .D(n9020), .Z(
        n8812) );
  HS65_LL_NOR4ABX2 U10184 ( .A(n9024), .B(n8993), .C(n14515), .D(n8812), .Z(
        n8271) );
  HS65_LL_NAND3X2 U10185 ( .A(n8828), .B(n8272), .C(n8271), .Z(n8307) );
  HS65_LL_IVX2 U10186 ( .A(n8273), .Z(n8841) );
  HS65_LL_AOI12X2 U10187 ( .A(n8300), .B(n12264), .C(n8841), .Z(n12273) );
  HS65_LL_NAND3X2 U10188 ( .A(n12273), .B(n8652), .C(n12279), .Z(n14505) );
  HS65_LL_NOR2X2 U10189 ( .A(n14526), .B(n8641), .Z(n15301) );
  HS65_LL_NOR3X1 U10190 ( .A(n15317), .B(n8275), .C(n8274), .Z(n8276) );
  HS65_LL_NAND3X2 U10191 ( .A(n8277), .B(n15301), .C(n8276), .Z(n9005) );
  HS65_LL_NOR2X2 U10192 ( .A(n12285), .B(n8987), .Z(n8278) );
  HS65_LL_NAND4ABX3 U10193 ( .A(n12278), .B(n9005), .C(n8278), .D(n15305), .Z(
        n8284) );
  HS65_LL_NAND2X2 U10194 ( .A(n12276), .B(n9025), .Z(n8661) );
  HS65_LL_NOR2X2 U10195 ( .A(n8279), .B(n8814), .Z(n12283) );
  HS65_LL_NAND2AX4 U10196 ( .A(n12283), .B(n15291), .Z(n14509) );
  HS65_LL_NOR2X2 U10197 ( .A(n8661), .B(n14509), .Z(n8813) );
  HS65_LL_NAND2X2 U10198 ( .A(sa13[1]), .B(n8281), .Z(n12274) );
  HS65_LL_OAI21X2 U10199 ( .A(sa13[7]), .B(n12274), .C(n12250), .Z(n14513) );
  HS65_LL_AOI12X2 U10200 ( .A(n8281), .B(n8663), .C(n8280), .Z(n8657) );
  HS65_LL_NOR3AX2 U10201 ( .A(n8657), .B(n8655), .C(n8282), .Z(n8283) );
  HS65_LL_NAND3X2 U10202 ( .A(n8283), .B(n8842), .C(n15278), .Z(n12288) );
  HS65_LL_NOR2X2 U10203 ( .A(n14513), .B(n12288), .Z(n8827) );
  HS65_LL_NAND4ABX3 U10204 ( .A(n14505), .B(n8284), .C(n8813), .D(n8827), .Z(
        n8306) );
  HS65_LL_NAND2X2 U10205 ( .A(n8286), .B(n8285), .Z(n8651) );
  HS65_LL_NAND2X2 U10206 ( .A(n8651), .B(n9007), .Z(n8646) );
  HS65_LL_NOR2X2 U10207 ( .A(n9006), .B(n8287), .Z(n8824) );
  HS65_LL_OAI112X1 U10208 ( .A(n8289), .B(n8288), .C(n8824), .D(n12239), .Z(
        n8294) );
  HS65_LL_NAND4ABX3 U10209 ( .A(n12283), .B(n8634), .C(n8992), .D(n9025), .Z(
        n8290) );
  HS65_LL_NOR4ABX2 U10210 ( .A(n8291), .B(n15305), .C(n8641), .D(n8290), .Z(
        n8292) );
  HS65_LL_NAND4ABX3 U10211 ( .A(n8646), .B(n8294), .C(n8293), .D(n8292), .Z(
        n8305) );
  HS65_LL_NAND2X2 U10212 ( .A(n8295), .B(n15304), .Z(n12244) );
  HS65_LL_NOR3X1 U10213 ( .A(n8996), .B(n8296), .C(n8995), .Z(n8983) );
  HS65_LL_OAI21X2 U10214 ( .A(n8988), .B(n9002), .C(n12266), .Z(n12253) );
  HS65_LL_NAND2X2 U10215 ( .A(n8298), .B(n8297), .Z(n8837) );
  HS65_LL_NAND4ABX3 U10216 ( .A(n8299), .B(n12253), .C(n8837), .D(n8805), .Z(
        n8665) );
  HS65_LL_NAND2X2 U10217 ( .A(n8300), .B(n8818), .Z(n8631) );
  HS65_LL_NAND3AX3 U10218 ( .A(n15293), .B(n8636), .C(n8631), .Z(n8301) );
  HS65_LL_NOR3X1 U10219 ( .A(n8983), .B(n8665), .C(n8301), .Z(n15311) );
  HS65_LL_NOR2X2 U10220 ( .A(n15281), .B(n8995), .Z(n8839) );
  HS65_LL_NOR4ABX2 U10221 ( .A(n15301), .B(n9024), .C(n8839), .D(n8302), .Z(
        n8303) );
  HS65_LL_NAND4ABX3 U10222 ( .A(n12244), .B(n8997), .C(n15311), .D(n8303), .Z(
        n8304) );
  HS65_LL_MX41X4 U10223 ( .D0(n8307), .S0(n15328), .D1(n8306), .S1(n15326), 
        .D2(n8305), .S2(n15324), .D3(n8304), .S3(n15322), .Z(n15277) );
  HS65_LL_MUXI21X2 U10224 ( .D0(n15648), .D1(n15649), .S0(n15277), .Z(n15579)
         );
  HS65_LL_IVX2 U10225 ( .A(n12307), .Z(n9047) );
  HS65_LL_NAND2X2 U10226 ( .A(n9047), .B(n15393), .Z(n8309) );
  HS65_LL_NAND4ABX3 U10227 ( .A(n12321), .B(n8309), .C(n15377), .D(n8308), .Z(
        n8310) );
  HS65_LL_NOR2X2 U10228 ( .A(n12308), .B(n9075), .Z(n9046) );
  HS65_LL_NAND4ABX3 U10229 ( .A(n8331), .B(n8310), .C(n9046), .D(n13032), .Z(
        n13043) );
  HS65_LL_NOR2X2 U10230 ( .A(n8312), .B(n8311), .Z(n8342) );
  HS65_LL_NAND4ABX3 U10231 ( .A(n8313), .B(n13043), .C(n8328), .D(n8342), .Z(
        n9043) );
  HS65_LL_NAND4ABX3 U10232 ( .A(n12301), .B(n9043), .C(n8315), .D(n8314), .Z(
        n8321) );
  HS65_LL_NOR2X2 U10233 ( .A(n8317), .B(n8316), .Z(n9054) );
  HS65_LL_NOR2AX3 U10234 ( .A(n12311), .B(n9054), .Z(n12337) );
  HS65_LL_NAND2X2 U10235 ( .A(n13019), .B(n8318), .Z(n12313) );
  HS65_LL_NAND2X2 U10236 ( .A(n8319), .B(n12313), .Z(n8337) );
  HS65_LL_NOR4ABX2 U10237 ( .A(n12337), .B(n15382), .C(n12316), .D(n8337), .Z(
        n9070) );
  HS65_LL_NAND4ABX3 U10238 ( .A(n8800), .B(n8321), .C(n9070), .D(n8320), .Z(
        n8351) );
  HS65_LL_NAND2X2 U10239 ( .A(n8322), .B(n8785), .Z(n15396) );
  HS65_LL_NOR2X2 U10240 ( .A(sa20[1]), .B(n15396), .Z(n9039) );
  HS65_LL_NOR2X2 U10241 ( .A(n9039), .B(n13031), .Z(n8332) );
  HS65_LL_NOR4ABX2 U10242 ( .A(n9062), .B(n8323), .C(n12308), .D(n13040), .Z(
        n8325) );
  HS65_LL_NOR4ABX2 U10243 ( .A(n8326), .B(n8325), .C(n8324), .D(n15418), .Z(
        n8327) );
  HS65_LL_NAND3X2 U10244 ( .A(n13038), .B(n8332), .C(n8327), .Z(n8350) );
  HS65_LL_NAND4ABX3 U10245 ( .A(n8329), .B(n12315), .C(n8328), .D(n9050), .Z(
        n8335) );
  HS65_LL_NOR2X2 U10246 ( .A(n9073), .B(n9054), .Z(n15385) );
  HS65_LL_NAND3X2 U10247 ( .A(sa20[5]), .B(sa20[0]), .C(n8330), .Z(n8345) );
  HS65_LL_NAND4ABX3 U10248 ( .A(n15384), .B(n8331), .C(n15385), .D(n8345), .Z(
        n8333) );
  HS65_LL_NAND4ABX3 U10249 ( .A(n8774), .B(n8333), .C(n8343), .D(n8332), .Z(
        n13021) );
  HS65_LL_NOR2X2 U10250 ( .A(n12307), .B(n13021), .Z(n8769) );
  HS65_LL_NOR4ABX2 U10251 ( .A(n8334), .B(n13036), .C(n8776), .D(n13040), .Z(
        n15404) );
  HS65_LL_NAND4ABX3 U10252 ( .A(n8336), .B(n8335), .C(n8769), .D(n15404), .Z(
        n8349) );
  HS65_LL_NOR2X2 U10253 ( .A(n8787), .B(n8337), .Z(n12293) );
  HS65_LL_NOR4ABX2 U10254 ( .A(n8340), .B(n15382), .C(n8339), .D(n8338), .Z(
        n8341) );
  HS65_LL_NAND3X2 U10255 ( .A(n8342), .B(n12293), .C(n8341), .Z(n8797) );
  HS65_LL_NAND4ABX3 U10256 ( .A(n13014), .B(n9039), .C(n8343), .D(n13025), .Z(
        n8347) );
  HS65_LL_NOR3X1 U10257 ( .A(sa20[6]), .B(n8784), .C(n8344), .Z(n8768) );
  HS65_LL_NOR4ABX2 U10258 ( .A(n8345), .B(n15377), .C(n8786), .D(n8768), .Z(
        n8346) );
  HS65_LL_NAND4ABX3 U10259 ( .A(n8797), .B(n8347), .C(n13047), .D(n8346), .Z(
        n8348) );
  HS65_LL_MX41X4 U10260 ( .D0(n8351), .S0(n13020), .D1(n8350), .S1(n15416), 
        .D2(n8349), .S2(n15408), .D3(n8348), .S3(n15400), .Z(n15421) );
  HS65_LLS_XOR3X2 U10261 ( .A(w2[19]), .B(n15579), .C(n15421), .Z(n8352) );
  HS65_LLS_XOR3X2 U10262 ( .A(n15630), .B(n14847), .C(n8352), .Z(n8353) );
  HS65_LL_MUX31X4 U10263 ( .D0(w2[19]), .D1(n15332), .D2(n8353), .S0(
        text_in_r[51]), .S1(n14808), .Z(N133) );
  HS65_LL_IVX2 U10264 ( .A(w0[26]), .Z(n15120) );
  HS65_LL_NAND2X2 U10265 ( .A(sa11[0]), .B(sa11[3]), .Z(n8355) );
  HS65_LL_IVX2 U10266 ( .A(n8355), .Z(n13591) );
  HS65_LL_NAND2X2 U10267 ( .A(sa11[5]), .B(n13591), .Z(n8383) );
  HS65_LL_NAND3X2 U10268 ( .A(sa11[1]), .B(sa11[6]), .C(sa11[7]), .Z(n11623)
         );
  HS65_LL_NOR2X2 U10269 ( .A(n8383), .B(n11623), .Z(n13602) );
  HS65_LL_NOR3X1 U10270 ( .A(sa11[1]), .B(sa11[6]), .C(sa11[7]), .Z(n11221) );
  HS65_LL_NOR3X1 U10271 ( .A(sa11[5]), .B(sa11[0]), .C(sa11[3]), .Z(n8371) );
  HS65_LL_NAND2X2 U10272 ( .A(n11221), .B(n8371), .Z(n13945) );
  HS65_LL_NOR2X2 U10273 ( .A(sa11[5]), .B(n8355), .Z(n8385) );
  HS65_LL_IVX2 U10274 ( .A(sa11[7]), .Z(n11215) );
  HS65_LL_NAND2X2 U10275 ( .A(sa11[6]), .B(n11215), .Z(n13579) );
  HS65_LL_NOR2X2 U10276 ( .A(sa11[1]), .B(n13579), .Z(n8377) );
  HS65_LL_NAND2X2 U10277 ( .A(n8385), .B(n8377), .Z(n11201) );
  HS65_LL_NAND2X2 U10278 ( .A(n13945), .B(n11201), .Z(n11619) );
  HS65_LL_NOR2X2 U10279 ( .A(n13602), .B(n11619), .Z(n12429) );
  HS65_LL_NOR2X2 U10280 ( .A(sa11[6]), .B(sa11[7]), .Z(n12976) );
  HS65_LL_NAND2X2 U10281 ( .A(sa11[1]), .B(n12976), .Z(n8366) );
  HS65_LL_IVX2 U10282 ( .A(sa11[3]), .Z(n12986) );
  HS65_LL_NOR2X2 U10283 ( .A(sa11[0]), .B(n12986), .Z(n11220) );
  HS65_LL_IVX2 U10284 ( .A(sa11[5]), .Z(n11624) );
  HS65_LL_NAND2X2 U10285 ( .A(n11220), .B(n11624), .Z(n11650) );
  HS65_LL_NOR2X2 U10286 ( .A(n8366), .B(n11650), .Z(n13942) );
  HS65_LL_NOR2X2 U10287 ( .A(sa11[0]), .B(sa11[3]), .Z(n12964) );
  HS65_LL_NAND2X2 U10288 ( .A(sa11[5]), .B(n12964), .Z(n8373) );
  HS65_LL_NOR2X2 U10289 ( .A(n8373), .B(n8366), .Z(n12981) );
  HS65_LL_IVX2 U10290 ( .A(sa11[1]), .Z(n8388) );
  HS65_LL_NOR2X2 U10291 ( .A(n8388), .B(n13579), .Z(n12963) );
  HS65_LL_IVX2 U10292 ( .A(n12963), .Z(n8381) );
  HS65_LL_NAND2X2 U10293 ( .A(sa11[5]), .B(n11220), .Z(n13578) );
  HS65_LL_NOR2X2 U10294 ( .A(n8381), .B(n13578), .Z(n11642) );
  HS65_LL_IVX2 U10295 ( .A(n11642), .Z(n8368) );
  HS65_LL_OR2X4 U10296 ( .A(n11623), .B(n11650), .Z(n11635) );
  HS65_LL_NAND2X2 U10297 ( .A(n8368), .B(n11635), .Z(n13971) );
  HS65_LL_NOR3X1 U10298 ( .A(n13942), .B(n12981), .C(n13971), .Z(n8354) );
  HS65_LL_NAND2X2 U10299 ( .A(sa11[0]), .B(n12986), .Z(n8357) );
  HS65_LL_NOR2X2 U10300 ( .A(sa11[5]), .B(n8357), .Z(n8378) );
  HS65_LL_NAND3X2 U10301 ( .A(sa11[6]), .B(sa11[7]), .C(n8378), .Z(n8394) );
  HS65_LL_NAND3X2 U10302 ( .A(n12429), .B(n8354), .C(n8394), .Z(n11216) );
  HS65_LL_NOR2X2 U10303 ( .A(sa11[6]), .B(n11215), .Z(n8379) );
  HS65_LL_NAND2X2 U10304 ( .A(n8379), .B(n8388), .Z(n8386) );
  HS65_LL_NOR2X2 U10305 ( .A(n8355), .B(n8386), .Z(n8527) );
  HS65_LL_IVX2 U10306 ( .A(n8366), .Z(n8372) );
  HS65_LL_NAND2X2 U10307 ( .A(sa11[5]), .B(n8372), .Z(n12985) );
  HS65_LL_NOR2X2 U10308 ( .A(n8355), .B(n12985), .Z(n13966) );
  HS65_LL_IVX2 U10309 ( .A(n8386), .Z(n8539) );
  HS65_LL_IVX2 U10310 ( .A(n11650), .Z(n12977) );
  HS65_LL_NAND2X2 U10311 ( .A(n8539), .B(n12977), .Z(n8533) );
  HS65_LL_IVX2 U10312 ( .A(n11221), .Z(n8367) );
  HS65_LL_NOR2X2 U10313 ( .A(n8367), .B(n13578), .Z(n13571) );
  HS65_LL_IVX2 U10314 ( .A(n13571), .Z(n8395) );
  HS65_LL_NAND2X2 U10315 ( .A(n8533), .B(n8395), .Z(n8530) );
  HS65_LL_IVX2 U10316 ( .A(n8530), .Z(n8356) );
  HS65_LL_IVX2 U10317 ( .A(n13579), .Z(n8358) );
  HS65_LL_NAND2X2 U10318 ( .A(n8358), .B(n12977), .Z(n12979) );
  HS65_LL_NAND4ABX3 U10319 ( .A(n8527), .B(n13966), .C(n8356), .D(n12979), .Z(
        n13948) );
  HS65_LL_NAND2X2 U10320 ( .A(sa11[1]), .B(n8379), .Z(n11649) );
  HS65_LL_NOR2X2 U10321 ( .A(n8373), .B(n11649), .Z(n13588) );
  HS65_LL_NOR2X2 U10322 ( .A(n8383), .B(n11649), .Z(n11206) );
  HS65_LL_IVX2 U10323 ( .A(n8385), .Z(n8521) );
  HS65_LL_NOR2X2 U10324 ( .A(n8521), .B(n8366), .Z(n11211) );
  HS65_LL_OR2X4 U10325 ( .A(n11206), .B(n11211), .Z(n13950) );
  HS65_LL_NOR2X2 U10326 ( .A(n13588), .B(n13950), .Z(n12970) );
  HS65_LL_IVX2 U10327 ( .A(n8383), .Z(n8362) );
  HS65_LL_NAND2X2 U10328 ( .A(n8362), .B(n11221), .Z(n12987) );
  HS65_LL_IVX2 U10329 ( .A(n8373), .Z(n8389) );
  HS65_LL_NAND2X2 U10330 ( .A(n8389), .B(n8539), .Z(n13965) );
  HS65_LL_IVX2 U10331 ( .A(n8357), .Z(n8361) );
  HS65_LL_NAND2X2 U10332 ( .A(n8361), .B(n11221), .Z(n11209) );
  HS65_LL_NOR2X2 U10333 ( .A(sa11[5]), .B(n11209), .Z(n12975) );
  HS65_LL_NAND2X2 U10334 ( .A(sa11[5]), .B(n8361), .Z(n11208) );
  HS65_LL_IVX2 U10335 ( .A(n11208), .Z(n8515) );
  HS65_LL_IVX2 U10336 ( .A(n8377), .Z(n11207) );
  HS65_LL_NOR2X2 U10337 ( .A(n8383), .B(n11207), .Z(n12417) );
  HS65_LL_AO12X4 U10338 ( .A(n8515), .B(n8358), .C(n12417), .Z(n8359) );
  HS65_LL_NOR4ABX2 U10339 ( .A(n12987), .B(n13965), .C(n12975), .D(n8359), .Z(
        n11654) );
  HS65_LL_NAND2X2 U10340 ( .A(n8515), .B(n8372), .Z(n8531) );
  HS65_LL_IVX2 U10341 ( .A(n8371), .Z(n8391) );
  HS65_LL_NOR2X2 U10342 ( .A(n11649), .B(n8391), .Z(n8363) );
  HS65_LL_IVX2 U10343 ( .A(n11209), .Z(n8376) );
  HS65_LL_NAND2X2 U10344 ( .A(sa11[5]), .B(n8376), .Z(n12403) );
  HS65_LL_NAND2X2 U10345 ( .A(n8371), .B(n8377), .Z(n12405) );
  HS65_LL_NAND2X2 U10346 ( .A(n12403), .B(n12405), .Z(n13970) );
  HS65_LL_NOR4ABX2 U10347 ( .A(n11654), .B(n8531), .C(n8363), .D(n13970), .Z(
        n8360) );
  HS65_LL_NAND4ABX3 U10348 ( .A(n11216), .B(n13948), .C(n12970), .D(n8360), 
        .Z(n8402) );
  HS65_LL_IVX2 U10349 ( .A(sa11[4]), .Z(n8397) );
  HS65_LL_NOR2X2 U10350 ( .A(sa11[2]), .B(n8397), .Z(n13972) );
  HS65_LL_NAND2X2 U10351 ( .A(n8361), .B(n8377), .Z(n8537) );
  HS65_LL_NOR2X2 U10352 ( .A(n11623), .B(n13578), .Z(n12997) );
  HS65_LL_NOR2X2 U10353 ( .A(n8381), .B(n11208), .Z(n12996) );
  HS65_LL_NAND2X2 U10354 ( .A(n8362), .B(n12963), .Z(n13958) );
  HS65_LL_NAND2X2 U10355 ( .A(n8378), .B(n8372), .Z(n13585) );
  HS65_LL_NAND2X2 U10356 ( .A(n13958), .B(n13585), .Z(n12956) );
  HS65_LL_NOR2X2 U10357 ( .A(n12996), .B(n12956), .Z(n12401) );
  HS65_LL_NOR2X2 U10358 ( .A(n8521), .B(n11623), .Z(n12412) );
  HS65_LL_NAND3X2 U10359 ( .A(sa11[6]), .B(sa11[7]), .C(n8388), .Z(n8520) );
  HS65_LL_NOR2X2 U10360 ( .A(n8520), .B(n13578), .Z(n12999) );
  HS65_LL_NOR2X2 U10361 ( .A(n12412), .B(n12999), .Z(n8374) );
  HS65_LL_IVX2 U10362 ( .A(n8363), .Z(n12423) );
  HS65_LL_NAND3X2 U10363 ( .A(n12401), .B(n8374), .C(n12423), .Z(n8364) );
  HS65_LL_NOR3AX2 U10364 ( .A(n8537), .B(n12997), .C(n8364), .Z(n13610) );
  HS65_LL_NAND2X2 U10365 ( .A(n12977), .B(n8377), .Z(n12422) );
  HS65_LL_NOR2X2 U10366 ( .A(n11208), .B(n11649), .Z(n12398) );
  HS65_LL_NOR4ABX2 U10367 ( .A(n8531), .B(n12422), .C(n12398), .D(n11206), .Z(
        n12394) );
  HS65_LL_NAND3X2 U10368 ( .A(sa11[5]), .B(n12963), .C(n12964), .Z(n11643) );
  HS65_LL_IVX2 U10369 ( .A(n8394), .Z(n12957) );
  HS65_LL_NAND2X2 U10370 ( .A(sa11[1]), .B(n12957), .Z(n8541) );
  HS65_LL_NAND2AX4 U10371 ( .A(n11619), .B(n8541), .Z(n13951) );
  HS65_LL_NOR4ABX2 U10372 ( .A(n12394), .B(n11643), .C(n8527), .D(n13951), .Z(
        n8365) );
  HS65_LL_NAND2X2 U10373 ( .A(n8378), .B(n12963), .Z(n8393) );
  HS65_LL_IVX2 U10374 ( .A(n8520), .Z(n8390) );
  HS65_LL_NAND2X2 U10375 ( .A(n8390), .B(n8371), .Z(n12955) );
  HS65_LL_NAND3X2 U10376 ( .A(n8365), .B(n8393), .C(n12955), .Z(n13975) );
  HS65_LL_NOR2X2 U10377 ( .A(n13588), .B(n13975), .Z(n12419) );
  HS65_LL_NOR2X2 U10378 ( .A(n8383), .B(n8520), .Z(n13599) );
  HS65_LL_NOR2X2 U10379 ( .A(sa11[3]), .B(n8366), .Z(n11626) );
  HS65_LL_NOR3X1 U10380 ( .A(sa11[6]), .B(n8388), .C(n11650), .Z(n12395) );
  HS65_LL_NOR3X1 U10381 ( .A(n13599), .B(n11626), .C(n12395), .Z(n8369) );
  HS65_LL_NAND2X2 U10382 ( .A(n12963), .B(n12977), .Z(n8524) );
  HS65_LL_NOR2X2 U10383 ( .A(n8367), .B(n8373), .Z(n13575) );
  HS65_LL_NOR3X1 U10384 ( .A(sa11[7]), .B(n8388), .C(n8521), .Z(n11628) );
  HS65_LL_NAND2X2 U10385 ( .A(n8515), .B(n8539), .Z(n13566) );
  HS65_LL_NAND2X2 U10386 ( .A(n8368), .B(n13566), .Z(n13604) );
  HS65_LL_NOR2X2 U10387 ( .A(n11628), .B(n13604), .Z(n12430) );
  HS65_LL_OR2X4 U10388 ( .A(n13578), .B(n8386), .Z(n13968) );
  HS65_LL_NAND2X2 U10389 ( .A(n12430), .B(n13968), .Z(n13983) );
  HS65_LL_NOR4ABX2 U10390 ( .A(n8369), .B(n8524), .C(n13575), .D(n13983), .Z(
        n8370) );
  HS65_LL_NAND3X2 U10391 ( .A(n13610), .B(n12419), .C(n8370), .Z(n8401) );
  HS65_LL_NOR2X2 U10392 ( .A(sa11[2]), .B(sa11[4]), .Z(n13961) );
  HS65_LL_IVX2 U10393 ( .A(n13575), .Z(n12954) );
  HS65_LL_NAND2X2 U10394 ( .A(n11643), .B(n12954), .Z(n12974) );
  HS65_LL_NOR2X2 U10395 ( .A(n8521), .B(n11649), .Z(n8516) );
  HS65_LL_IVX2 U10396 ( .A(n13566), .Z(n13967) );
  HS65_LL_NOR2X2 U10397 ( .A(n8516), .B(n13967), .Z(n12958) );
  HS65_LL_NOR2X2 U10398 ( .A(n8381), .B(n8391), .Z(n13598) );
  HS65_LL_AOI12X2 U10399 ( .A(n8386), .B(n11207), .C(n8391), .Z(n12988) );
  HS65_LL_NAND2X2 U10400 ( .A(n8372), .B(n8371), .Z(n13943) );
  HS65_LL_NAND2X2 U10401 ( .A(n11221), .B(n12977), .Z(n13593) );
  HS65_LL_NAND2X2 U10402 ( .A(n13943), .B(n13593), .Z(n13568) );
  HS65_LL_NOR2X2 U10403 ( .A(n8373), .B(n11623), .Z(n8382) );
  HS65_LL_IVX2 U10404 ( .A(n8524), .Z(n11634) );
  HS65_LL_NOR2X2 U10405 ( .A(n8382), .B(n11634), .Z(n11195) );
  HS65_LL_NAND4ABX3 U10406 ( .A(n12988), .B(n13568), .C(n8374), .D(n11195), 
        .Z(n8375) );
  HS65_LL_NOR3X1 U10407 ( .A(n8376), .B(n13598), .C(n8375), .Z(n12393) );
  HS65_LL_NOR2X2 U10408 ( .A(sa11[5]), .B(n8537), .Z(n13583) );
  HS65_LL_NAND2X2 U10409 ( .A(n8390), .B(n12977), .Z(n12410) );
  HS65_LL_IVX2 U10410 ( .A(n11649), .Z(n13590) );
  HS65_LL_NAND2X2 U10411 ( .A(n8378), .B(n13590), .Z(n11203) );
  HS65_LL_NAND2X2 U10412 ( .A(n12410), .B(n11203), .Z(n11224) );
  HS65_LL_NAND2X2 U10413 ( .A(n8389), .B(n8377), .Z(n11636) );
  HS65_LL_NAND2X2 U10414 ( .A(n11221), .B(n8385), .Z(n11646) );
  HS65_LL_NAND2X2 U10415 ( .A(n11636), .B(n11646), .Z(n11223) );
  HS65_LL_NOR3X1 U10416 ( .A(n13583), .B(n11224), .C(n11223), .Z(n13969) );
  HS65_LL_NAND2X2 U10417 ( .A(n8379), .B(n8378), .Z(n8517) );
  HS65_LL_NOR2X2 U10418 ( .A(sa11[1]), .B(n8517), .Z(n11644) );
  HS65_LL_NOR4ABX2 U10419 ( .A(n12393), .B(n13969), .C(n11644), .D(n11211), 
        .Z(n8380) );
  HS65_LL_NAND4ABX3 U10420 ( .A(n11216), .B(n12974), .C(n12958), .D(n8380), 
        .Z(n8400) );
  HS65_LL_IVX2 U10421 ( .A(sa11[2]), .Z(n8398) );
  HS65_LL_NOR2X2 U10422 ( .A(sa11[4]), .B(n8398), .Z(n13614) );
  HS65_LL_IVX2 U10423 ( .A(n12987), .Z(n12960) );
  HS65_LL_NOR2X2 U10424 ( .A(n8521), .B(n8381), .Z(n12416) );
  HS65_LL_NOR2X2 U10425 ( .A(n12960), .B(n12416), .Z(n13577) );
  HS65_LL_NOR2X2 U10426 ( .A(n8520), .B(n11208), .Z(n12990) );
  HS65_LL_NOR2X2 U10427 ( .A(n12990), .B(n8382), .Z(n12400) );
  HS65_LL_NOR2X2 U10428 ( .A(n8383), .B(n8386), .Z(n13003) );
  HS65_LL_IVX2 U10429 ( .A(n8531), .Z(n13605) );
  HS65_LL_NOR3X1 U10430 ( .A(n11644), .B(n13003), .C(n13605), .Z(n8384) );
  HS65_LL_NAND3X2 U10431 ( .A(n13577), .B(n12400), .C(n8384), .Z(n11219) );
  HS65_LL_NAND2X2 U10432 ( .A(n8385), .B(n8539), .Z(n11202) );
  HS65_LL_NAND2AX4 U10433 ( .A(n12412), .B(n11202), .Z(n12425) );
  HS65_LL_NOR2X2 U10434 ( .A(n11649), .B(n13578), .Z(n12962) );
  HS65_LL_NOR2X2 U10435 ( .A(n8386), .B(n8391), .Z(n11637) );
  HS65_LL_NOR2X2 U10436 ( .A(n12962), .B(n11637), .Z(n12406) );
  HS65_LL_NAND3X2 U10437 ( .A(n12406), .B(n8541), .C(n13958), .Z(n8387) );
  HS65_LL_NOR3X1 U10438 ( .A(n12395), .B(n12425), .C(n8387), .Z(n8551) );
  HS65_LL_NAND3X2 U10439 ( .A(sa11[6]), .B(n12977), .C(n8388), .Z(n11639) );
  HS65_LL_NAND2X2 U10440 ( .A(n8551), .B(n11639), .Z(n12973) );
  HS65_LL_NOR2AX3 U10441 ( .A(n11220), .B(n12985), .Z(n11200) );
  HS65_LL_IVX2 U10442 ( .A(n13945), .Z(n12989) );
  HS65_LL_NOR2X2 U10443 ( .A(n12417), .B(n12989), .Z(n12959) );
  HS65_LL_NAND2X2 U10444 ( .A(n12959), .B(n8533), .Z(n13963) );
  HS65_LL_NAND2X2 U10445 ( .A(n8390), .B(n8389), .Z(n12418) );
  HS65_LL_IVX2 U10446 ( .A(n8516), .Z(n11645) );
  HS65_LL_NAND2X2 U10447 ( .A(n12418), .B(n11645), .Z(n11656) );
  HS65_LL_NOR3X1 U10448 ( .A(n11200), .B(n13963), .C(n11656), .Z(n8392) );
  HS65_LL_NOR2X2 U10449 ( .A(n11623), .B(n8391), .Z(n13941) );
  HS65_LL_IVX2 U10450 ( .A(n13941), .Z(n11630) );
  HS65_LL_NAND3X2 U10451 ( .A(n8392), .B(n12403), .C(n11630), .Z(n13612) );
  HS65_LL_IVX2 U10452 ( .A(n8393), .Z(n11625) );
  HS65_LL_NOR2X2 U10453 ( .A(sa11[1]), .B(n8394), .Z(n13576) );
  HS65_LL_NOR3X1 U10454 ( .A(n12997), .B(n11625), .C(n13576), .Z(n8526) );
  HS65_LL_NAND3X2 U10455 ( .A(n8526), .B(n13943), .C(n8395), .Z(n11652) );
  HS65_LL_NOR2X2 U10456 ( .A(n13612), .B(n11652), .Z(n12984) );
  HS65_LL_IVX2 U10457 ( .A(n13588), .Z(n8536) );
  HS65_LL_NOR4ABX2 U10458 ( .A(n11636), .B(n8536), .C(n11642), .D(n13602), .Z(
        n8396) );
  HS65_LL_NAND4ABX3 U10459 ( .A(n11219), .B(n12973), .C(n12984), .D(n8396), 
        .Z(n8399) );
  HS65_LL_NOR2X2 U10460 ( .A(n8398), .B(n8397), .Z(n13981) );
  HS65_LL_MX41X4 U10461 ( .D0(n8402), .S0(n13972), .D1(n8401), .S1(n13961), 
        .D2(n8400), .S2(n13614), .D3(n8399), .S3(n13981), .Z(n15259) );
  HS65_LL_IVX2 U10462 ( .A(sa00[7]), .Z(n12864) );
  HS65_LL_NAND2X2 U10463 ( .A(sa00[6]), .B(n12864), .Z(n11154) );
  HS65_LL_IVX2 U10464 ( .A(n11154), .Z(n11156) );
  HS65_LL_NAND2X2 U10465 ( .A(sa00[1]), .B(n11156), .Z(n12872) );
  HS65_LL_IVX2 U10466 ( .A(sa00[3]), .Z(n11177) );
  HS65_LL_NOR2X2 U10467 ( .A(sa00[0]), .B(n11177), .Z(n11159) );
  HS65_LL_NAND2X2 U10468 ( .A(sa00[5]), .B(n11159), .Z(n11183) );
  HS65_LL_NOR2X2 U10469 ( .A(n12872), .B(n11183), .Z(n12568) );
  HS65_LL_IVX2 U10470 ( .A(sa00[1]), .Z(n13693) );
  HS65_LL_NAND2X2 U10471 ( .A(sa00[7]), .B(n13693), .Z(n11184) );
  HS65_LL_NOR2X2 U10472 ( .A(sa00[6]), .B(n11184), .Z(n11160) );
  HS65_LL_IVX2 U10473 ( .A(n11160), .Z(n8421) );
  HS65_LL_IVX2 U10474 ( .A(sa00[5]), .Z(n8427) );
  HS65_LL_NAND3X2 U10475 ( .A(sa00[3]), .B(sa00[0]), .C(n8427), .Z(n12578) );
  HS65_LL_NOR2X2 U10476 ( .A(n8421), .B(n12578), .Z(n11161) );
  HS65_LL_IVX2 U10477 ( .A(sa00[6]), .Z(n13692) );
  HS65_LL_NAND3X2 U10478 ( .A(sa00[7]), .B(sa00[1]), .C(n13692), .Z(n11150) );
  HS65_LL_NOR2X2 U10479 ( .A(n11183), .B(n11150), .Z(n11175) );
  HS65_LL_NOR2X2 U10480 ( .A(n11161), .B(n11175), .Z(n12877) );
  HS65_LL_NAND3X2 U10481 ( .A(sa00[1]), .B(sa00[7]), .C(sa00[6]), .Z(n11188)
         );
  HS65_LL_NOR2X2 U10482 ( .A(n11188), .B(n12578), .Z(n11174) );
  HS65_LL_NAND2X2 U10483 ( .A(n11159), .B(n8427), .Z(n8428) );
  HS65_LL_NOR2X2 U10484 ( .A(n8428), .B(n11150), .Z(n13467) );
  HS65_LL_NOR2X2 U10485 ( .A(n11174), .B(n13467), .Z(n13670) );
  HS65_LL_NOR2X2 U10486 ( .A(sa00[3]), .B(sa00[0]), .Z(n12869) );
  HS65_LL_NAND2X2 U10487 ( .A(n12869), .B(n8427), .Z(n12572) );
  HS65_LL_IVX2 U10488 ( .A(n12572), .Z(n12586) );
  HS65_LL_NAND2X2 U10489 ( .A(n11160), .B(n12586), .Z(n13487) );
  HS65_LL_IVX2 U10490 ( .A(n8428), .Z(n13702) );
  HS65_LL_NOR3X1 U10491 ( .A(sa00[7]), .B(sa00[6]), .C(n13693), .Z(n8417) );
  HS65_LL_NAND2X2 U10492 ( .A(n13702), .B(n8417), .Z(n13986) );
  HS65_LL_NAND3X2 U10493 ( .A(sa00[5]), .B(sa00[3]), .C(sa00[0]), .Z(n8418) );
  HS65_LL_NOR2X2 U10494 ( .A(n12872), .B(n8418), .Z(n13695) );
  HS65_LL_IVX2 U10495 ( .A(sa00[0]), .Z(n8408) );
  HS65_LL_NOR2X2 U10496 ( .A(sa00[3]), .B(n8408), .Z(n8404) );
  HS65_LL_NAND2X2 U10497 ( .A(n8404), .B(n8427), .Z(n13665) );
  HS65_LL_NOR2X2 U10498 ( .A(n11188), .B(n13665), .Z(n14095) );
  HS65_LL_NOR4ABX2 U10499 ( .A(n13487), .B(n13986), .C(n13695), .D(n14095), 
        .Z(n8403) );
  HS65_LL_NAND3X2 U10500 ( .A(n12877), .B(n13670), .C(n8403), .Z(n14132) );
  HS65_LL_NAND2X2 U10501 ( .A(sa00[5]), .B(n12869), .Z(n11155) );
  HS65_LL_NOR3X1 U10502 ( .A(n11154), .B(n11155), .C(sa00[1]), .Z(n13479) );
  HS65_LL_IVX2 U10503 ( .A(n13479), .Z(n12544) );
  HS65_LL_NOR2X2 U10504 ( .A(n13692), .B(n8428), .Z(n13668) );
  HS65_LL_NAND2X2 U10505 ( .A(n13668), .B(n13693), .Z(n13490) );
  HS65_LL_NOR2X2 U10506 ( .A(n11155), .B(n11150), .Z(n14094) );
  HS65_LL_NOR2X2 U10507 ( .A(n8418), .B(n11188), .Z(n13677) );
  HS65_LL_NOR4ABX2 U10508 ( .A(n12544), .B(n13490), .C(n14094), .D(n13677), 
        .Z(n8407) );
  HS65_LL_NOR2X2 U10509 ( .A(n8421), .B(n13665), .Z(n13481) );
  HS65_LL_IVX2 U10510 ( .A(n8404), .Z(n11180) );
  HS65_LL_NOR2X2 U10511 ( .A(n8427), .B(n11180), .Z(n8424) );
  HS65_LL_NAND2X2 U10512 ( .A(n8424), .B(n8417), .Z(n11171) );
  HS65_LL_IVX2 U10513 ( .A(n8418), .Z(n8413) );
  HS65_LL_NAND2X2 U10514 ( .A(n8413), .B(n11160), .Z(n12893) );
  HS65_LL_NAND2X2 U10515 ( .A(n11171), .B(n12893), .Z(n8410) );
  HS65_LL_NOR2X2 U10516 ( .A(n11155), .B(n11188), .Z(n13683) );
  HS65_LL_NAND3X2 U10517 ( .A(sa00[7]), .B(sa00[6]), .C(n13693), .Z(n14115) );
  HS65_LL_IVX2 U10518 ( .A(n8424), .Z(n11187) );
  HS65_LL_NOR2X2 U10519 ( .A(n14115), .B(n11187), .Z(n12583) );
  HS65_LL_NOR2X2 U10520 ( .A(n13683), .B(n12583), .Z(n12558) );
  HS65_LL_NOR2X2 U10521 ( .A(n12872), .B(n12578), .Z(n13672) );
  HS65_LL_NAND3X2 U10522 ( .A(n13693), .B(n12864), .C(n13692), .Z(n12554) );
  HS65_LL_NOR2X2 U10523 ( .A(n12554), .B(n8418), .Z(n12874) );
  HS65_LL_NOR2X2 U10524 ( .A(n13672), .B(n12874), .Z(n8405) );
  HS65_LL_NAND4ABX3 U10525 ( .A(n13481), .B(n8410), .C(n12558), .D(n8405), .Z(
        n11190) );
  HS65_LL_IVX2 U10526 ( .A(n11159), .Z(n12555) );
  HS65_LL_NAND2X2 U10527 ( .A(sa00[5]), .B(n8417), .Z(n11176) );
  HS65_LL_NOR2X2 U10528 ( .A(n11188), .B(n12572), .Z(n12867) );
  HS65_LL_IVX2 U10529 ( .A(n12867), .Z(n12884) );
  HS65_LL_IVX2 U10530 ( .A(n12554), .Z(n8426) );
  HS65_LL_NAND2X2 U10531 ( .A(n8426), .B(n8424), .Z(n12579) );
  HS65_LL_OAI112X1 U10532 ( .A(n12555), .B(n11176), .C(n12884), .D(n12579), 
        .Z(n14120) );
  HS65_LL_NOR2X2 U10533 ( .A(sa00[1]), .B(n11154), .Z(n12585) );
  HS65_LL_NAND2X2 U10534 ( .A(n12585), .B(n8413), .Z(n12894) );
  HS65_LL_NAND2X2 U10535 ( .A(n8426), .B(n12586), .Z(n13684) );
  HS65_LL_NAND2X2 U10536 ( .A(n12894), .B(n13684), .Z(n12870) );
  HS65_LL_NOR2X2 U10537 ( .A(n14115), .B(n11155), .Z(n11178) );
  HS65_LL_NOR2X2 U10538 ( .A(n11150), .B(n12578), .Z(n13497) );
  HS65_LL_NOR2X2 U10539 ( .A(n11178), .B(n13497), .Z(n14127) );
  HS65_LL_NAND2X2 U10540 ( .A(n13702), .B(n11160), .Z(n13997) );
  HS65_LL_NAND4ABX3 U10541 ( .A(n14120), .B(n12870), .C(n14127), .D(n13997), 
        .Z(n12549) );
  HS65_LL_NOR2X2 U10542 ( .A(n14115), .B(n13665), .Z(n14105) );
  HS65_LL_NOR2X2 U10543 ( .A(n11188), .B(n11183), .Z(n13661) );
  HS65_LL_NOR2X2 U10544 ( .A(n12872), .B(n13665), .Z(n13478) );
  HS65_LL_NOR3X1 U10545 ( .A(n14105), .B(n13661), .C(n13478), .Z(n12883) );
  HS65_LL_NAND2X2 U10546 ( .A(n8417), .B(n12586), .Z(n14114) );
  HS65_LL_IVX2 U10547 ( .A(n11183), .Z(n13699) );
  HS65_LL_NAND2X2 U10548 ( .A(n8426), .B(n13699), .Z(n12587) );
  HS65_LL_NAND3X2 U10549 ( .A(n12883), .B(n14114), .C(n12587), .Z(n13471) );
  HS65_LL_NOR3X1 U10550 ( .A(n11190), .B(n12549), .C(n13471), .Z(n8406) );
  HS65_LL_NAND4ABX3 U10551 ( .A(n12568), .B(n14132), .C(n8407), .D(n8406), .Z(
        n8436) );
  HS65_LL_NAND2X2 U10552 ( .A(sa00[2]), .B(sa00[4]), .Z(n14134) );
  HS65_LL_IVX2 U10553 ( .A(n14134), .Z(n13709) );
  HS65_LL_IVX2 U10554 ( .A(n12578), .Z(n12865) );
  HS65_LL_AOI12X2 U10555 ( .A(n12865), .B(n12585), .C(n13478), .Z(n12557) );
  HS65_LL_NAND3AX3 U10556 ( .A(n11161), .B(n12557), .C(n13684), .Z(n11181) );
  HS65_LL_NOR2X2 U10557 ( .A(n14115), .B(n12572), .Z(n14104) );
  HS65_LL_NOR2X2 U10558 ( .A(n14095), .B(n14104), .Z(n12875) );
  HS65_LL_NOR2X2 U10559 ( .A(n12872), .B(n11155), .Z(n12584) );
  HS65_LL_IVX2 U10560 ( .A(n12585), .Z(n14108) );
  HS65_LL_NOR2X2 U10561 ( .A(n14108), .B(n8428), .Z(n12891) );
  HS65_LL_NOR3X1 U10562 ( .A(n8427), .B(n8408), .C(n11150), .Z(n13701) );
  HS65_LL_NOR3X1 U10563 ( .A(n12584), .B(n12891), .C(n13701), .Z(n8409) );
  HS65_LL_NAND4ABX3 U10564 ( .A(n8410), .B(n11181), .C(n12875), .D(n8409), .Z(
        n14010) );
  HS65_LL_NOR2X2 U10565 ( .A(n8428), .B(n12872), .Z(n11169) );
  HS65_LL_NOR2X2 U10566 ( .A(n11183), .B(n8421), .Z(n14003) );
  HS65_LL_NOR2X2 U10567 ( .A(n11169), .B(n14003), .Z(n12882) );
  HS65_LL_NOR2X2 U10568 ( .A(n12554), .B(n11155), .Z(n12564) );
  HS65_LL_IVX2 U10569 ( .A(n13986), .Z(n8411) );
  HS65_LL_NOR2X2 U10570 ( .A(n12564), .B(n8411), .Z(n12550) );
  HS65_LL_NAND4ABX3 U10571 ( .A(n14094), .B(n13467), .C(n12882), .D(n12550), 
        .Z(n8415) );
  HS65_LL_NOR3X1 U10572 ( .A(sa00[7]), .B(n13693), .C(n12578), .Z(n8412) );
  HS65_LL_IVX2 U10573 ( .A(n12568), .Z(n12588) );
  HS65_LL_NOR2X2 U10574 ( .A(n11180), .B(n8421), .Z(n11170) );
  HS65_LL_NAND2X2 U10575 ( .A(sa00[5]), .B(n11170), .Z(n12871) );
  HS65_LL_NAND2X2 U10576 ( .A(n12588), .B(n12871), .Z(n14002) );
  HS65_LL_NOR2X2 U10577 ( .A(n8412), .B(n14002), .Z(n13994) );
  HS65_LL_NOR2X2 U10578 ( .A(n14108), .B(n11180), .Z(n11163) );
  HS65_LL_NAND2AX4 U10579 ( .A(n11150), .B(n12586), .Z(n13996) );
  HS65_LL_IVX2 U10580 ( .A(n11174), .Z(n8429) );
  HS65_LL_NAND2X2 U10581 ( .A(n13996), .B(n8429), .Z(n13682) );
  HS65_LL_NOR2X2 U10582 ( .A(n12872), .B(n11187), .Z(n14097) );
  HS65_LL_IVX2 U10583 ( .A(n13665), .Z(n8422) );
  HS65_LL_NAND2X2 U10584 ( .A(n8417), .B(n8422), .Z(n13488) );
  HS65_LL_IVX2 U10585 ( .A(n13488), .Z(n13998) );
  HS65_LL_NOR3X1 U10586 ( .A(n14097), .B(n13998), .C(n13695), .Z(n12560) );
  HS65_LL_NOR2X2 U10587 ( .A(n14115), .B(n11183), .Z(n12561) );
  HS65_LL_NOR2X2 U10588 ( .A(n12561), .B(n13661), .Z(n12896) );
  HS65_LL_NAND4ABX3 U10589 ( .A(n11163), .B(n13682), .C(n12560), .D(n12896), 
        .Z(n13474) );
  HS65_LL_IVX2 U10590 ( .A(n13474), .Z(n8414) );
  HS65_LL_IVX2 U10591 ( .A(n14115), .Z(n11152) );
  HS65_LL_NAND2X2 U10592 ( .A(n11152), .B(n8413), .Z(n13685) );
  HS65_LL_NAND2X2 U10593 ( .A(n8414), .B(n13685), .Z(n12553) );
  HS65_LL_AOI12X2 U10594 ( .A(n12869), .B(n8417), .C(n12553), .Z(n13483) );
  HS65_LL_NAND4ABX3 U10595 ( .A(n14010), .B(n8415), .C(n13994), .D(n13483), 
        .Z(n8435) );
  HS65_LL_NOR2X2 U10596 ( .A(sa00[2]), .B(sa00[4]), .Z(n14130) );
  HS65_LL_NOR2AX3 U10597 ( .A(n12893), .B(n11169), .Z(n12545) );
  HS65_LL_IVX2 U10598 ( .A(n8417), .Z(n8419) );
  HS65_LL_NOR2X2 U10599 ( .A(n8418), .B(n8419), .Z(n14004) );
  HS65_LL_NAND2X2 U10600 ( .A(n13997), .B(n12587), .Z(n14122) );
  HS65_LL_NOR3X1 U10601 ( .A(n11161), .B(n14004), .C(n14122), .Z(n8416) );
  HS65_LL_IVX2 U10602 ( .A(n12891), .Z(n13694) );
  HS65_LL_NAND3X2 U10603 ( .A(n12545), .B(n8416), .C(n13694), .Z(n13992) );
  HS65_LL_IVX2 U10604 ( .A(n11171), .Z(n13697) );
  HS65_LL_OAI21X2 U10605 ( .A(n14108), .B(n12572), .C(n12579), .Z(n14007) );
  HS65_LL_NAND2X2 U10606 ( .A(n8417), .B(n12865), .Z(n14013) );
  HS65_LL_NOR2X2 U10607 ( .A(n8418), .B(n11150), .Z(n14012) );
  HS65_LL_NOR3AX2 U10608 ( .A(n14013), .B(n14094), .C(n14012), .Z(n12885) );
  HS65_LL_NAND4ABX3 U10609 ( .A(n13697), .B(n14007), .C(n12885), .D(n13996), 
        .Z(n8425) );
  HS65_LL_NOR2X2 U10610 ( .A(n8428), .B(n11188), .Z(n14000) );
  HS65_LL_NOR2X2 U10611 ( .A(n11155), .B(n8419), .Z(n12582) );
  HS65_LL_AOI12X2 U10612 ( .A(n12865), .B(n12585), .C(n12582), .Z(n13499) );
  HS65_LL_NAND2X2 U10613 ( .A(n13499), .B(n13684), .Z(n13477) );
  HS65_LL_NOR2X2 U10614 ( .A(n14095), .B(n13477), .Z(n14016) );
  HS65_LL_NAND4ABX3 U10615 ( .A(n14105), .B(n14000), .C(n13986), .D(n14016), 
        .Z(n8420) );
  HS65_LL_NOR3X1 U10616 ( .A(n12568), .B(n13677), .C(n8420), .Z(n11185) );
  HS65_LL_NOR2X2 U10617 ( .A(n11155), .B(n8421), .Z(n14001) );
  HS65_LL_NAND2X2 U10618 ( .A(n8426), .B(n8422), .Z(n13662) );
  HS65_LL_NAND4ABX3 U10619 ( .A(n14001), .B(n12874), .C(n13662), .D(n12894), 
        .Z(n8423) );
  HS65_LL_AOI12X2 U10620 ( .A(n11156), .B(n8424), .C(n8423), .Z(n13469) );
  HS65_LL_NAND4ABX3 U10621 ( .A(n13992), .B(n8425), .C(n11185), .D(n13469), 
        .Z(n8434) );
  HS65_LL_IVX2 U10622 ( .A(sa00[2]), .Z(n8432) );
  HS65_LL_NAND2X2 U10623 ( .A(sa00[4]), .B(n8432), .Z(n14125) );
  HS65_LL_IVX2 U10624 ( .A(n14125), .Z(n14008) );
  HS65_LL_NAND2X2 U10625 ( .A(n8426), .B(n12865), .Z(n11173) );
  HS65_LL_AND2X4 U10626 ( .A(n11173), .B(n12544), .Z(n11151) );
  HS65_LL_NOR2X2 U10627 ( .A(n13665), .B(n11150), .Z(n14096) );
  HS65_LL_NOR2X2 U10628 ( .A(n8428), .B(n14115), .Z(n11164) );
  HS65_LL_NOR2X2 U10629 ( .A(n14096), .B(n11164), .Z(n13681) );
  HS65_LL_NAND2X2 U10630 ( .A(n8427), .B(n11163), .Z(n11162) );
  HS65_LL_NAND3X2 U10631 ( .A(n11151), .B(n13681), .C(n11162), .Z(n14006) );
  HS65_LL_NOR2AX3 U10632 ( .A(n13487), .B(n12561), .Z(n11167) );
  HS65_LL_NAND2X2 U10633 ( .A(n11167), .B(n14114), .Z(n13999) );
  HS65_LL_NOR2X2 U10634 ( .A(n13683), .B(n14007), .Z(n13482) );
  HS65_LL_NOR2X2 U10635 ( .A(n8428), .B(n12554), .Z(n12548) );
  HS65_LL_NOR2X2 U10636 ( .A(n12872), .B(n12572), .Z(n12546) );
  HS65_LL_NOR4ABX2 U10637 ( .A(n13482), .B(n13662), .C(n12548), .D(n12546), 
        .Z(n8430) );
  HS65_LL_NAND4ABX3 U10638 ( .A(n11169), .B(n13999), .C(n8430), .D(n8429), .Z(
        n13705) );
  HS65_LL_NOR2X2 U10639 ( .A(n12564), .B(n13497), .Z(n13663) );
  HS65_LL_NOR4ABX2 U10640 ( .A(n13663), .B(n14013), .C(n11170), .D(n12584), 
        .Z(n8431) );
  HS65_LL_NAND4ABX3 U10641 ( .A(n14006), .B(n13705), .C(n11185), .D(n8431), 
        .Z(n8433) );
  HS65_LL_NOR2X2 U10642 ( .A(sa00[4]), .B(n8432), .Z(n14137) );
  HS65_LL_MX41X4 U10643 ( .D0(n8436), .S0(n13709), .D1(n8435), .S1(n14130), 
        .D2(n8434), .S2(n14008), .D3(n8433), .S3(n14137), .Z(n15552) );
  HS65_LL_IVX2 U10644 ( .A(sa33[1]), .Z(n11266) );
  HS65_LL_NOR2X2 U10645 ( .A(n11266), .B(sa33[7]), .Z(n8458) );
  HS65_LL_IVX2 U10646 ( .A(n8458), .Z(n13559) );
  HS65_LL_NOR2X2 U10647 ( .A(sa33[6]), .B(n13559), .Z(n13517) );
  HS65_LL_IVX2 U10648 ( .A(sa33[0]), .Z(n8437) );
  HS65_LL_NAND2X2 U10649 ( .A(sa33[5]), .B(n8437), .Z(n14040) );
  HS65_LL_NOR2X2 U10650 ( .A(sa33[3]), .B(n14040), .Z(n11231) );
  HS65_LL_NAND2X2 U10651 ( .A(n13517), .B(n11231), .Z(n13544) );
  HS65_LL_NAND2X2 U10652 ( .A(sa33[5]), .B(sa33[0]), .Z(n11293) );
  HS65_LL_IVX2 U10653 ( .A(n11293), .Z(n12596) );
  HS65_LL_NAND3X2 U10654 ( .A(n13517), .B(sa33[3]), .C(n12596), .Z(n11289) );
  HS65_LL_NOR2X2 U10655 ( .A(sa33[5]), .B(n8437), .Z(n13554) );
  HS65_LL_NAND2X2 U10656 ( .A(sa33[3]), .B(n13554), .Z(n8440) );
  HS65_LL_NOR2X2 U10657 ( .A(n13559), .B(n8440), .Z(n13533) );
  HS65_LL_NAND2X2 U10658 ( .A(sa33[6]), .B(n13533), .Z(n13626) );
  HS65_LL_NAND3X2 U10659 ( .A(n13544), .B(n11289), .C(n13626), .Z(n13525) );
  HS65_LL_IVX2 U10660 ( .A(n13517), .Z(n8455) );
  HS65_LL_IVX2 U10661 ( .A(sa33[3]), .Z(n8459) );
  HS65_LL_NAND2X2 U10662 ( .A(n12596), .B(n8459), .Z(n11258) );
  HS65_LL_NOR2X2 U10663 ( .A(n8455), .B(n11258), .Z(n11717) );
  HS65_LL_IVX2 U10664 ( .A(n13554), .Z(n12611) );
  HS65_LL_NOR2X2 U10665 ( .A(sa33[3]), .B(n12611), .Z(n8469) );
  HS65_LL_IVX2 U10666 ( .A(sa33[6]), .Z(n8439) );
  HS65_LL_NAND3X2 U10667 ( .A(sa33[7]), .B(n8469), .C(n8439), .Z(n8461) );
  HS65_LL_NOR2X2 U10668 ( .A(sa33[1]), .B(n8461), .Z(n12621) );
  HS65_LL_IVX2 U10669 ( .A(n11231), .Z(n13558) );
  HS65_LL_NAND3X2 U10670 ( .A(sa33[6]), .B(sa33[1]), .C(sa33[7]), .Z(n8468) );
  HS65_LL_NOR2X2 U10671 ( .A(n13558), .B(n8468), .Z(n13640) );
  HS65_LL_NOR3X1 U10672 ( .A(n11717), .B(n12621), .C(n13640), .Z(n11259) );
  HS65_LL_NAND2X2 U10673 ( .A(sa33[3]), .B(n12596), .Z(n11297) );
  HS65_LL_NAND3X2 U10674 ( .A(sa33[6]), .B(sa33[7]), .C(n11266), .Z(n11721) );
  HS65_LL_NOR2X2 U10675 ( .A(n11297), .B(n11721), .Z(n13639) );
  HS65_LL_NAND2X2 U10676 ( .A(sa33[6]), .B(n8458), .Z(n11243) );
  HS65_LL_IVX2 U10677 ( .A(n14040), .Z(n8463) );
  HS65_LL_NAND2X2 U10678 ( .A(sa33[3]), .B(n8463), .Z(n11722) );
  HS65_LL_NOR2X2 U10679 ( .A(n11243), .B(n11722), .Z(n13650) );
  HS65_LL_NOR2X2 U10680 ( .A(n13639), .B(n13650), .Z(n13549) );
  HS65_LL_IVX2 U10681 ( .A(n8469), .Z(n8445) );
  HS65_LL_NOR2X2 U10682 ( .A(sa33[1]), .B(n8439), .Z(n14036) );
  HS65_LL_IVX2 U10683 ( .A(n14036), .Z(n14057) );
  HS65_LL_NOR2X2 U10684 ( .A(n14057), .B(sa33[7]), .Z(n11270) );
  HS65_LL_IVX2 U10685 ( .A(n11270), .Z(n11287) );
  HS65_LL_NOR2X2 U10686 ( .A(n8445), .B(n11287), .Z(n14044) );
  HS65_LL_NOR2X2 U10687 ( .A(sa33[5]), .B(sa33[0]), .Z(n13518) );
  HS65_LL_NAND2X2 U10688 ( .A(sa33[3]), .B(n13518), .Z(n14058) );
  HS65_LL_NOR2X2 U10689 ( .A(n14058), .B(n11243), .Z(n11276) );
  HS65_LL_NOR3X1 U10690 ( .A(sa33[6]), .B(sa33[1]), .C(sa33[7]), .Z(n11237) );
  HS65_LL_IVX2 U10691 ( .A(n14058), .Z(n11275) );
  HS65_LL_NAND2X2 U10692 ( .A(n11237), .B(n11275), .Z(n13621) );
  HS65_LL_IVX2 U10693 ( .A(n11258), .Z(n8444) );
  HS65_LL_NAND3X2 U10694 ( .A(n8439), .B(n11266), .C(sa33[7]), .Z(n8442) );
  HS65_LL_IVX2 U10695 ( .A(n8442), .Z(n13555) );
  HS65_LL_NAND2X2 U10696 ( .A(n8444), .B(n13555), .Z(n11727) );
  HS65_LL_NAND2X2 U10697 ( .A(n13621), .B(n11727), .Z(n8449) );
  HS65_LL_NOR3X1 U10698 ( .A(n14044), .B(n11276), .C(n8449), .Z(n8438) );
  HS65_LL_NAND3X2 U10699 ( .A(n11259), .B(n13549), .C(n8438), .Z(n11256) );
  HS65_LL_NAND3X2 U10700 ( .A(sa33[1]), .B(sa33[7]), .C(n8439), .Z(n14039) );
  HS65_LL_NOR2X2 U10701 ( .A(n8445), .B(n14039), .Z(n11285) );
  HS65_LL_NOR2X2 U10702 ( .A(n11258), .B(n11243), .Z(n14030) );
  HS65_LL_NOR2X2 U10703 ( .A(n11285), .B(n14030), .Z(n11235) );
  HS65_LL_NOR2X2 U10704 ( .A(n8468), .B(n11297), .Z(n13630) );
  HS65_LL_NOR2X2 U10705 ( .A(n8440), .B(n8442), .Z(n11291) );
  HS65_LL_NOR2X2 U10706 ( .A(n13630), .B(n11291), .Z(n13637) );
  HS65_LL_NAND2X2 U10707 ( .A(n11237), .B(n8444), .Z(n11720) );
  HS65_LL_IVX2 U10708 ( .A(n8440), .Z(n14035) );
  HS65_LL_NAND2X2 U10709 ( .A(n13517), .B(n14035), .Z(n13632) );
  HS65_LL_NAND2X2 U10710 ( .A(n11231), .B(n11237), .Z(n11708) );
  HS65_LL_NAND2X2 U10711 ( .A(n13632), .B(n11708), .Z(n11728) );
  HS65_LL_NOR2X2 U10712 ( .A(n8440), .B(n11721), .Z(n11278) );
  HS65_LL_NOR2X2 U10713 ( .A(n11258), .B(n8468), .Z(n13537) );
  HS65_LL_NOR2X2 U10714 ( .A(n11278), .B(n13537), .Z(n11260) );
  HS65_LL_NOR2X2 U10715 ( .A(n8442), .B(n11297), .Z(n11290) );
  HS65_LL_NOR2X2 U10716 ( .A(n11297), .B(n11287), .Z(n11712) );
  HS65_LL_NOR2X2 U10717 ( .A(n11290), .B(n11712), .Z(n14029) );
  HS65_LL_IVX2 U10718 ( .A(n11237), .Z(n8450) );
  HS65_LL_NOR2X2 U10719 ( .A(n8440), .B(n8450), .Z(n13551) );
  HS65_LL_NAND2X2 U10720 ( .A(n13518), .B(n8459), .Z(n11725) );
  HS65_LL_NOR2X2 U10721 ( .A(n8468), .B(n11725), .Z(n14062) );
  HS65_LL_NOR2X2 U10722 ( .A(n13551), .B(n14062), .Z(n8447) );
  HS65_LL_NAND3X2 U10723 ( .A(n11260), .B(n14029), .C(n8447), .Z(n8441) );
  HS65_LL_NOR4ABX2 U10724 ( .A(n13637), .B(n11720), .C(n11728), .D(n8441), .Z(
        n13521) );
  HS65_LL_NOR2X2 U10725 ( .A(n8445), .B(n8468), .Z(n13629) );
  HS65_LL_NOR2X2 U10726 ( .A(n13558), .B(n14039), .Z(n11715) );
  HS65_LL_NOR2X2 U10727 ( .A(n13629), .B(n11715), .Z(n8453) );
  HS65_LL_NAND3X2 U10728 ( .A(n11235), .B(n13521), .C(n8453), .Z(n8473) );
  HS65_LL_NOR2X2 U10729 ( .A(n14058), .B(n8442), .Z(n11283) );
  HS65_LL_IVX2 U10730 ( .A(n11722), .Z(n8467) );
  HS65_LL_IVX2 U10731 ( .A(n14039), .Z(n8460) );
  HS65_LL_NAND2X2 U10732 ( .A(n8467), .B(n8460), .Z(n13619) );
  HS65_LL_IVX2 U10733 ( .A(n13619), .Z(n14048) );
  HS65_LL_NOR2X2 U10734 ( .A(n11283), .B(n14048), .Z(n8472) );
  HS65_LL_IVX2 U10735 ( .A(n11725), .Z(n11239) );
  HS65_LL_NAND2X2 U10736 ( .A(n8460), .B(n11239), .Z(n12607) );
  HS65_LL_OAI21X2 U10737 ( .A(n11722), .B(n11721), .C(n12607), .Z(n11246) );
  HS65_LL_NAND2X2 U10738 ( .A(n13517), .B(n8469), .Z(n12617) );
  HS65_LL_NAND2X2 U10739 ( .A(n13517), .B(n11239), .Z(n8448) );
  HS65_LL_NAND2X2 U10740 ( .A(n13555), .B(n11239), .Z(n11279) );
  HS65_LL_NAND3X2 U10741 ( .A(n12617), .B(n8448), .C(n11279), .Z(n8443) );
  HS65_LL_NOR3AX2 U10742 ( .A(n8472), .B(n11246), .C(n8443), .Z(n11301) );
  HS65_LL_NAND2X2 U10743 ( .A(n8444), .B(n8460), .Z(n13511) );
  HS65_LL_NAND2X2 U10744 ( .A(n8444), .B(n11270), .Z(n13631) );
  HS65_LL_NOR2X2 U10745 ( .A(n8445), .B(n11721), .Z(n12606) );
  HS65_LL_NOR2X2 U10746 ( .A(n11721), .B(n11725), .Z(n14054) );
  HS65_LL_NOR4ABX2 U10747 ( .A(n13511), .B(n13631), .C(n12606), .D(n14054), 
        .Z(n8446) );
  HS65_LL_NAND4ABX3 U10748 ( .A(n11256), .B(n8473), .C(n11301), .D(n8446), .Z(
        n8479) );
  HS65_LL_NOR2AX3 U10749 ( .A(sa33[2]), .B(sa33[4]), .Z(n14075) );
  HS65_LL_IVX2 U10750 ( .A(n8447), .Z(n14027) );
  HS65_LL_NAND2AX4 U10751 ( .A(n8468), .B(n14035), .Z(n13641) );
  HS65_LL_NAND2X2 U10752 ( .A(n13619), .B(n13641), .Z(n8457) );
  HS65_LL_NOR2X2 U10753 ( .A(n14027), .B(n8457), .Z(n12615) );
  HS65_LL_IVX2 U10754 ( .A(n8448), .Z(n13541) );
  HS65_LL_NOR2X2 U10755 ( .A(n13541), .B(n8449), .Z(n12610) );
  HS65_LL_NAND2X2 U10756 ( .A(n14035), .B(n11270), .Z(n13528) );
  HS65_LL_NOR2X2 U10757 ( .A(n14058), .B(n8468), .Z(n13526) );
  HS65_LL_NAND2X2 U10758 ( .A(sa33[7]), .B(n8467), .Z(n14031) );
  HS65_LL_NOR3X1 U10759 ( .A(sa33[6]), .B(sa33[1]), .C(n14031), .Z(n12629) );
  HS65_LL_IVX2 U10760 ( .A(n13525), .Z(n14060) );
  HS65_LL_NOR2X2 U10761 ( .A(n13558), .B(n11721), .Z(n8466) );
  HS65_LL_NOR2X2 U10762 ( .A(n14058), .B(n11721), .Z(n13529) );
  HS65_LL_IVX2 U10763 ( .A(n13631), .Z(n11244) );
  HS65_LL_NAND2X2 U10764 ( .A(n11231), .B(n13555), .Z(n8465) );
  HS65_LL_OAI21X2 U10765 ( .A(n11721), .B(n11258), .C(n8465), .Z(n11252) );
  HS65_LL_NOR2X2 U10766 ( .A(n11244), .B(n11252), .Z(n14059) );
  HS65_LL_NOR2X2 U10767 ( .A(n8450), .B(n11297), .Z(n14047) );
  HS65_LL_NOR2X2 U10768 ( .A(n14044), .B(n14047), .Z(n12613) );
  HS65_LL_NAND3X2 U10769 ( .A(n13637), .B(n14059), .C(n12613), .Z(n8451) );
  HS65_LL_NOR3X1 U10770 ( .A(n8466), .B(n13529), .C(n8451), .Z(n13654) );
  HS65_LL_IVX2 U10771 ( .A(n11720), .Z(n11288) );
  HS65_LL_NOR2X2 U10772 ( .A(n11288), .B(n11283), .Z(n11251) );
  HS65_LL_NAND3X2 U10773 ( .A(n14060), .B(n13654), .C(n11251), .Z(n8452) );
  HS65_LL_NOR3X1 U10774 ( .A(n14030), .B(n12629), .C(n8452), .Z(n11234) );
  HS65_LL_OAI112X1 U10775 ( .A(n11297), .B(n14057), .C(n8453), .D(n11234), .Z(
        n8454) );
  HS65_LL_NOR4ABX2 U10776 ( .A(n12610), .B(n13528), .C(n13526), .D(n8454), .Z(
        n8477) );
  HS65_LL_NAND2X2 U10777 ( .A(sa33[4]), .B(sa33[2]), .Z(n14079) );
  HS65_LL_NOR2X2 U10778 ( .A(sa33[4]), .B(sa33[2]), .Z(n13657) );
  HS65_LL_NOR2X2 U10779 ( .A(n11291), .B(n13629), .Z(n14046) );
  HS65_LL_IVX2 U10780 ( .A(n11279), .Z(n11723) );
  HS65_LL_NOR2X2 U10781 ( .A(n11297), .B(n11243), .Z(n14034) );
  HS65_LL_NAND2X2 U10782 ( .A(n11275), .B(n8460), .Z(n13506) );
  HS65_LL_NOR2X2 U10783 ( .A(n8455), .B(n8459), .Z(n12625) );
  HS65_LL_NAND2X2 U10784 ( .A(n13518), .B(n12625), .Z(n14028) );
  HS65_LL_NAND2X2 U10785 ( .A(n13506), .B(n14028), .Z(n13648) );
  HS65_LL_NOR3X1 U10786 ( .A(n11723), .B(n14034), .C(n13648), .Z(n8456) );
  HS65_LL_NAND3AX3 U10787 ( .A(n8457), .B(n14046), .C(n8456), .Z(n14069) );
  HS65_LL_IVX2 U10788 ( .A(n11717), .Z(n11292) );
  HS65_LL_IVX2 U10789 ( .A(n14062), .Z(n11248) );
  HS65_LL_NAND2X2 U10790 ( .A(n11292), .B(n11248), .Z(n13532) );
  HS65_LL_AOI12X2 U10791 ( .A(n8458), .B(n11239), .C(n11278), .Z(n13508) );
  HS65_LL_NOR2X2 U10792 ( .A(n11722), .B(n11287), .Z(n13516) );
  HS65_LL_NOR2X2 U10793 ( .A(n13639), .B(n13516), .Z(n12612) );
  HS65_LL_NOR2X2 U10794 ( .A(n11276), .B(n11283), .Z(n11272) );
  HS65_LL_NAND2X2 U10795 ( .A(n8463), .B(n11237), .Z(n12608) );
  HS65_LL_NOR3X1 U10796 ( .A(sa33[0]), .B(n8459), .C(n8468), .Z(n13647) );
  HS65_LL_NAND2X2 U10797 ( .A(n11237), .B(n8469), .Z(n12600) );
  HS65_LL_NAND2X2 U10798 ( .A(n13631), .B(n12600), .Z(n11713) );
  HS65_LL_NOR4ABX2 U10799 ( .A(n11272), .B(n12608), .C(n13647), .D(n11713), 
        .Z(n8462) );
  HS65_LL_NAND2X2 U10800 ( .A(n14035), .B(n8460), .Z(n13548) );
  HS65_LL_NAND3X2 U10801 ( .A(n8462), .B(n8461), .C(n13548), .Z(n13625) );
  HS65_LL_IVX2 U10802 ( .A(n14047), .Z(n11714) );
  HS65_LL_NAND2X2 U10803 ( .A(n8463), .B(n12625), .Z(n11249) );
  HS65_LL_NAND2X2 U10804 ( .A(n11714), .B(n11249), .Z(n13519) );
  HS65_LL_NOR4ABX2 U10805 ( .A(n12612), .B(n11720), .C(n13625), .D(n13519), 
        .Z(n8464) );
  HS65_LL_NAND4ABX3 U10806 ( .A(n14069), .B(n13532), .C(n13508), .D(n8464), 
        .Z(n8475) );
  HS65_LL_NOR2AX3 U10807 ( .A(sa33[4]), .B(sa33[2]), .Z(n14067) );
  HS65_LL_IVX2 U10808 ( .A(n8465), .Z(n13543) );
  HS65_LL_IVX2 U10809 ( .A(n8466), .Z(n13618) );
  HS65_LL_NAND2X2 U10810 ( .A(n13618), .B(n13548), .Z(n13515) );
  HS65_LL_NOR2X2 U10811 ( .A(n13526), .B(n13515), .Z(n13507) );
  HS65_LL_NAND2X2 U10812 ( .A(n11237), .B(n8467), .Z(n13527) );
  HS65_LL_IVX2 U10813 ( .A(n12607), .Z(n11716) );
  HS65_LL_IVX2 U10814 ( .A(n12617), .Z(n14050) );
  HS65_LL_NOR2X2 U10815 ( .A(n14050), .B(n12629), .Z(n11281) );
  HS65_LL_NOR2X2 U10816 ( .A(n8468), .B(n11722), .Z(n11247) );
  HS65_LL_NOR2X2 U10817 ( .A(n12606), .B(n11247), .Z(n11703) );
  HS65_LL_IVX2 U10818 ( .A(n13516), .Z(n11282) );
  HS65_LL_IVX2 U10819 ( .A(n11243), .Z(n11240) );
  HS65_LL_NAND2X2 U10820 ( .A(n8469), .B(n11240), .Z(n11702) );
  HS65_LL_NAND2X2 U10821 ( .A(n11282), .B(n11702), .Z(n12598) );
  HS65_LL_NAND2X2 U10822 ( .A(n13621), .B(n13511), .Z(n11241) );
  HS65_LL_NOR3X1 U10823 ( .A(n11276), .B(n12598), .C(n11241), .Z(n8470) );
  HS65_LL_NAND3X2 U10824 ( .A(n11281), .B(n11703), .C(n8470), .Z(n14066) );
  HS65_LL_NOR4ABX2 U10825 ( .A(n13507), .B(n13527), .C(n11716), .D(n14066), 
        .Z(n8471) );
  HS65_LL_NAND4ABX3 U10826 ( .A(n13543), .B(n8473), .C(n8472), .D(n8471), .Z(
        n8474) );
  HS65_LL_AOI22X1 U10827 ( .A(n13657), .B(n8475), .C(n14067), .D(n8474), .Z(
        n8476) );
  HS65_LL_CBI4I1X3 U10828 ( .A(n12615), .B(n8477), .C(n14079), .D(n8476), .Z(
        n8478) );
  HS65_LL_CBI4I6X2 U10829 ( .A(n13525), .B(n8479), .C(n14075), .D(n8478), .Z(
        n14819) );
  HS65_LL_NOR2X2 U10830 ( .A(sa22[2]), .B(sa22[4]), .Z(n12945) );
  HS65_LL_IVX2 U10831 ( .A(sa22[3]), .Z(n10128) );
  HS65_LL_NAND2X2 U10832 ( .A(sa22[0]), .B(n10128), .Z(n10134) );
  HS65_LL_NOR2X2 U10833 ( .A(sa22[5]), .B(n10134), .Z(n8502) );
  HS65_LL_IVX2 U10834 ( .A(n8502), .Z(n11675) );
  HS65_LL_IVX2 U10835 ( .A(sa22[1]), .Z(n11667) );
  HS65_LL_NAND2X2 U10836 ( .A(sa22[6]), .B(sa22[7]), .Z(n11674) );
  HS65_LL_NOR2X2 U10837 ( .A(n11667), .B(n11674), .Z(n8489) );
  HS65_LL_IVX2 U10838 ( .A(n8489), .Z(n8496) );
  HS65_LL_NOR2X2 U10839 ( .A(n11675), .B(n8496), .Z(n11321) );
  HS65_LL_IVX2 U10840 ( .A(sa22[6]), .Z(n8480) );
  HS65_LL_NAND2X2 U10841 ( .A(sa22[7]), .B(n8480), .Z(n10101) );
  HS65_LL_NOR2X2 U10842 ( .A(sa22[1]), .B(n10101), .Z(n10108) );
  HS65_LL_NAND2X2 U10843 ( .A(sa22[3]), .B(sa22[0]), .Z(n11324) );
  HS65_LL_NOR2X2 U10844 ( .A(sa22[5]), .B(n11324), .Z(n10087) );
  HS65_LL_NAND2X2 U10845 ( .A(n10108), .B(n10087), .Z(n11661) );
  HS65_LL_NAND2AX4 U10846 ( .A(n11321), .B(n11661), .Z(n12927) );
  HS65_LL_NOR2X2 U10847 ( .A(sa22[0]), .B(n10128), .Z(n10131) );
  HS65_LL_IVX2 U10848 ( .A(sa22[5]), .Z(n10129) );
  HS65_LL_NAND2X2 U10849 ( .A(n10131), .B(n10129), .Z(n10111) );
  HS65_LL_NOR3X1 U10850 ( .A(sa22[6]), .B(n11667), .C(n10111), .Z(n12451) );
  HS65_LL_NAND2X2 U10851 ( .A(sa22[5]), .B(n10131), .Z(n8495) );
  HS65_LL_IVX2 U10852 ( .A(n10101), .Z(n8498) );
  HS65_LL_NAND2X2 U10853 ( .A(sa22[1]), .B(n8498), .Z(n11323) );
  HS65_LL_NOR2X2 U10854 ( .A(n8495), .B(n11323), .Z(n12913) );
  HS65_LL_IVX2 U10855 ( .A(n10108), .Z(n10119) );
  HS65_LL_NOR2X2 U10856 ( .A(sa22[3]), .B(sa22[0]), .Z(n12930) );
  HS65_LL_NAND2X2 U10857 ( .A(n12930), .B(n10129), .Z(n10112) );
  HS65_LL_NOR2X2 U10858 ( .A(n10119), .B(n10112), .Z(n10135) );
  HS65_LL_NOR2X2 U10859 ( .A(n12913), .B(n10135), .Z(n11692) );
  HS65_LL_NAND2X2 U10860 ( .A(n10087), .B(n8489), .Z(n11665) );
  HS65_LL_NOR2X2 U10861 ( .A(n10129), .B(n11324), .Z(n12923) );
  HS65_LL_NOR2X2 U10862 ( .A(n8480), .B(sa22[7]), .Z(n8482) );
  HS65_LL_IVX2 U10863 ( .A(n8482), .Z(n10118) );
  HS65_LL_NOR2X2 U10864 ( .A(n11667), .B(n10118), .Z(n12929) );
  HS65_LL_NAND2X2 U10865 ( .A(n12923), .B(n12929), .Z(n12448) );
  HS65_LL_NAND3X2 U10866 ( .A(n11692), .B(n11665), .C(n12448), .Z(n8481) );
  HS65_LL_NOR3X1 U10867 ( .A(n12927), .B(n12451), .C(n8481), .Z(n12920) );
  HS65_LL_NOR2X2 U10868 ( .A(sa22[6]), .B(sa22[7]), .Z(n12500) );
  HS65_LL_NAND2X2 U10869 ( .A(n12500), .B(n11667), .Z(n10133) );
  HS65_LL_NAND2X2 U10870 ( .A(sa22[5]), .B(n12930), .Z(n10117) );
  HS65_LL_NOR2X2 U10871 ( .A(n10133), .B(n10117), .Z(n12526) );
  HS65_LL_NOR2X2 U10872 ( .A(n10119), .B(n10111), .Z(n11343) );
  HS65_LL_IVX2 U10873 ( .A(n10087), .Z(n8490) );
  HS65_LL_NOR2X2 U10874 ( .A(n11323), .B(n8490), .Z(n11743) );
  HS65_LL_IVX2 U10875 ( .A(n10111), .Z(n11309) );
  HS65_LL_NAND2X2 U10876 ( .A(n8489), .B(n11309), .Z(n10122) );
  HS65_LL_IVX2 U10877 ( .A(n10122), .Z(n10099) );
  HS65_LL_OR3X4 U10878 ( .A(n11343), .B(n11743), .C(n10099), .Z(n8504) );
  HS65_LL_AOI112X2 U10879 ( .A(n8502), .B(n8498), .C(n12526), .D(n8504), .Z(
        n8483) );
  HS65_LL_NAND2X2 U10880 ( .A(n8482), .B(n11667), .Z(n10091) );
  HS65_LL_NOR2X2 U10881 ( .A(n10134), .B(n10091), .Z(n10092) );
  HS65_LL_NAND2X2 U10882 ( .A(sa22[5]), .B(n10092), .Z(n12477) );
  HS65_LL_IVX2 U10883 ( .A(n8495), .Z(n11745) );
  HS65_LL_IVX2 U10884 ( .A(n10133), .Z(n12922) );
  HS65_LL_NAND2X2 U10885 ( .A(n11745), .B(n12922), .Z(n10116) );
  HS65_LL_NOR2X2 U10886 ( .A(n8495), .B(n11674), .Z(n12936) );
  HS65_LL_NAND2X2 U10887 ( .A(sa22[1]), .B(n12936), .Z(n12449) );
  HS65_LL_NAND2X2 U10888 ( .A(n10116), .B(n12449), .Z(n10095) );
  HS65_LL_NAND2X2 U10889 ( .A(n11309), .B(n12929), .Z(n10121) );
  HS65_LL_NAND2X2 U10890 ( .A(n8502), .B(n12922), .Z(n12515) );
  HS65_LL_NAND2X2 U10891 ( .A(n10121), .B(n12515), .Z(n11749) );
  HS65_LL_NOR4ABX2 U10892 ( .A(n8483), .B(n12477), .C(n10095), .D(n11749), .Z(
        n12464) );
  HS65_LL_IVX2 U10893 ( .A(n12923), .Z(n10124) );
  HS65_LL_IVX2 U10894 ( .A(n11674), .Z(n10088) );
  HS65_LL_NAND2X2 U10895 ( .A(n10088), .B(n11667), .Z(n8485) );
  HS65_LL_NOR2X2 U10896 ( .A(n10124), .B(n8485), .Z(n12441) );
  HS65_LL_IVX2 U10897 ( .A(n10112), .Z(n10107) );
  HS65_LL_NAND2X2 U10898 ( .A(n10107), .B(n12929), .Z(n12467) );
  HS65_LL_IVX2 U10899 ( .A(n12467), .Z(n11318) );
  HS65_LL_NOR2X2 U10900 ( .A(n12441), .B(n11318), .Z(n12521) );
  HS65_LL_NAND2X2 U10901 ( .A(sa22[1]), .B(n12500), .Z(n10110) );
  HS65_LL_NOR2X2 U10902 ( .A(n10112), .B(n10110), .Z(n11747) );
  HS65_LL_NOR2X2 U10903 ( .A(n8495), .B(n10110), .Z(n11689) );
  HS65_LL_IVX2 U10904 ( .A(n10091), .Z(n11340) );
  HS65_LL_NAND2X2 U10905 ( .A(n11745), .B(n11340), .Z(n11322) );
  HS65_LL_NAND2X2 U10906 ( .A(n12923), .B(n12922), .Z(n11669) );
  HS65_LL_NAND2X2 U10907 ( .A(n11322), .B(n11669), .Z(n12487) );
  HS65_LL_NOR3X1 U10908 ( .A(n11747), .B(n11689), .C(n12487), .Z(n10109) );
  HS65_LL_NOR2X2 U10909 ( .A(n10129), .B(n10134), .Z(n8488) );
  HS65_LL_IVX2 U10910 ( .A(n8488), .Z(n10100) );
  HS65_LL_NOR3X1 U10911 ( .A(sa22[6]), .B(sa22[7]), .C(n10100), .Z(n11737) );
  HS65_LL_NOR2X2 U10912 ( .A(n10112), .B(n8496), .Z(n11334) );
  HS65_LL_IVX2 U10913 ( .A(n8485), .Z(n11746) );
  HS65_LL_NAND2X2 U10914 ( .A(n10087), .B(n11746), .Z(n12911) );
  HS65_LL_IVX2 U10915 ( .A(n12911), .Z(n12446) );
  HS65_LL_OR2X4 U10916 ( .A(n11334), .B(n12446), .Z(n12917) );
  HS65_LL_NOR4ABX2 U10917 ( .A(n12521), .B(n10109), .C(n11737), .D(n12917), 
        .Z(n8484) );
  HS65_LL_NAND3X2 U10918 ( .A(n12920), .B(n12464), .C(n8484), .Z(n8514) );
  HS65_LL_IVX2 U10919 ( .A(n11665), .Z(n12472) );
  HS65_LL_NOR2X2 U10920 ( .A(n8490), .B(n10133), .Z(n11308) );
  HS65_LL_NOR2X2 U10921 ( .A(n11334), .B(n11308), .Z(n8491) );
  HS65_LL_IVX2 U10922 ( .A(n12913), .Z(n11679) );
  HS65_LL_NAND2X2 U10923 ( .A(n8491), .B(n11679), .Z(n11666) );
  HS65_LL_NOR2X2 U10924 ( .A(n12472), .B(n11666), .Z(n12495) );
  HS65_LL_NOR3X1 U10925 ( .A(sa22[1]), .B(n10101), .C(n10100), .Z(n12530) );
  HS65_LL_IVX2 U10926 ( .A(n12441), .Z(n11331) );
  HS65_LL_NAND2X2 U10927 ( .A(n11309), .B(n12922), .Z(n12527) );
  HS65_LL_NAND2X2 U10928 ( .A(n11331), .B(n12527), .Z(n12511) );
  HS65_LL_NOR2X2 U10929 ( .A(n12530), .B(n12511), .Z(n8497) );
  HS65_LL_NOR2X2 U10930 ( .A(n11323), .B(n10117), .Z(n11761) );
  HS65_LL_NOR2X2 U10931 ( .A(n11321), .B(n11761), .Z(n8493) );
  HS65_LL_NOR2X2 U10932 ( .A(n10133), .B(n10100), .Z(n11744) );
  HS65_LL_NOR2X2 U10933 ( .A(n11343), .B(n11744), .Z(n11684) );
  HS65_LL_NOR2X2 U10934 ( .A(n10119), .B(n10117), .Z(n12462) );
  HS65_LL_NOR2X2 U10935 ( .A(n8485), .B(n10100), .Z(n12504) );
  HS65_LL_NOR2X2 U10936 ( .A(n12462), .B(n12504), .Z(n11680) );
  HS65_LL_NOR2X2 U10937 ( .A(n10117), .B(n8485), .Z(n10127) );
  HS65_LL_NOR3X1 U10938 ( .A(sa22[1]), .B(n11674), .C(n10111), .Z(n11307) );
  HS65_LL_NOR3X1 U10939 ( .A(n10092), .B(n10127), .C(n11307), .Z(n8486) );
  HS65_LL_IVX2 U10940 ( .A(n11669), .Z(n10096) );
  HS65_LL_NAND2X2 U10941 ( .A(n8489), .B(n12923), .Z(n10120) );
  HS65_LL_NAND2X2 U10942 ( .A(n11661), .B(n10120), .Z(n12513) );
  HS65_LL_NOR4ABX2 U10943 ( .A(n11680), .B(n8486), .C(n10096), .D(n12513), .Z(
        n12457) );
  HS65_LL_IVX2 U10944 ( .A(n12929), .Z(n8494) );
  HS65_LL_NOR2X2 U10945 ( .A(n8494), .B(n10100), .Z(n10098) );
  HS65_LL_NOR2X2 U10946 ( .A(n8490), .B(n8494), .Z(n12492) );
  HS65_LL_NOR2X2 U10947 ( .A(n10110), .B(n10117), .Z(n12505) );
  HS65_LL_NOR2X2 U10948 ( .A(n10110), .B(n10124), .Z(n12524) );
  HS65_LL_NOR3X1 U10949 ( .A(n12492), .B(n12505), .C(n12524), .Z(n12915) );
  HS65_LL_NAND2X2 U10950 ( .A(n11745), .B(n10108), .Z(n12501) );
  HS65_LL_NAND2X2 U10951 ( .A(n12915), .B(n12501), .Z(n10104) );
  HS65_LL_NOR4ABX2 U10952 ( .A(n11684), .B(n12457), .C(n10098), .D(n10104), 
        .Z(n11695) );
  HS65_LL_OAI112X1 U10953 ( .A(n11324), .B(n10091), .C(n8493), .D(n11695), .Z(
        n8487) );
  HS65_LL_NOR4ABX2 U10954 ( .A(n8497), .B(n10122), .C(n11747), .D(n8487), .Z(
        n8512) );
  HS65_LL_NAND2X2 U10955 ( .A(sa22[2]), .B(sa22[4]), .Z(n11339) );
  HS65_LL_NOR2X2 U10956 ( .A(n11323), .B(n11675), .Z(n12485) );
  HS65_LL_NOR2X2 U10957 ( .A(n10098), .B(n12485), .Z(n10125) );
  HS65_LL_NAND2X2 U10958 ( .A(n8489), .B(n8488), .Z(n12533) );
  HS65_LL_NAND2X2 U10959 ( .A(n12911), .B(n12533), .Z(n10093) );
  HS65_LL_NOR2X2 U10960 ( .A(n10124), .B(n10091), .Z(n12460) );
  HS65_LL_NOR3X1 U10961 ( .A(n11667), .B(n8490), .C(sa22[7]), .Z(n11335) );
  HS65_LL_NOR2AX3 U10962 ( .A(n11335), .B(sa22[6]), .Z(n11751) );
  HS65_LL_NOR2X2 U10963 ( .A(n12460), .B(n11751), .Z(n11663) );
  HS65_LL_NOR2X2 U10964 ( .A(n10119), .B(n10124), .Z(n11310) );
  HS65_LL_NOR2AX3 U10965 ( .A(n8491), .B(n11310), .Z(n12939) );
  HS65_LL_NAND4ABX3 U10966 ( .A(n10093), .B(n12513), .C(n11663), .D(n12939), 
        .Z(n8492) );
  HS65_LL_NOR3X1 U10967 ( .A(n12526), .B(n11744), .C(n8492), .Z(n12509) );
  HS65_LL_NAND3X2 U10968 ( .A(n10125), .B(n12509), .C(n8493), .Z(n8510) );
  HS65_LL_NOR2X2 U10969 ( .A(n11323), .B(n10100), .Z(n12469) );
  HS65_LL_IVX2 U10970 ( .A(n12915), .Z(n12535) );
  HS65_LL_NAND2X2 U10971 ( .A(n8502), .B(n11746), .Z(n12473) );
  HS65_LL_NAND2X2 U10972 ( .A(n8502), .B(n11340), .Z(n12458) );
  HS65_LL_NAND2X2 U10973 ( .A(n10121), .B(n12458), .Z(n12908) );
  HS65_LL_NOR2X2 U10974 ( .A(n8495), .B(n8494), .Z(n12498) );
  HS65_LL_NOR2X2 U10975 ( .A(n10110), .B(n10100), .Z(n12453) );
  HS65_LL_OR2X4 U10976 ( .A(n12498), .B(n12453), .Z(n12512) );
  HS65_LL_NOR2X2 U10977 ( .A(n8496), .B(n10117), .Z(n12440) );
  HS65_LL_AOI12X2 U10978 ( .A(n8502), .B(n10108), .C(n12440), .Z(n10090) );
  HS65_LL_NAND4ABX3 U10979 ( .A(n12908), .B(n12512), .C(n8497), .D(n10090), 
        .Z(n11664) );
  HS65_LL_IVX2 U10980 ( .A(n10110), .Z(n10130) );
  HS65_LL_NAND2X2 U10981 ( .A(n8502), .B(n10130), .Z(n10123) );
  HS65_LL_NOR2AX3 U10982 ( .A(n10123), .B(n12913), .Z(n12925) );
  HS65_LL_CBI4I6X2 U10983 ( .A(n8498), .B(n10130), .C(n10107), .D(n11343), .Z(
        n8500) );
  HS65_LL_NAND2X2 U10984 ( .A(n11745), .B(n11746), .Z(n8499) );
  HS65_LL_NAND3X2 U10985 ( .A(n12925), .B(n8500), .C(n8499), .Z(n11325) );
  HS65_LL_NOR4ABX2 U10986 ( .A(n12477), .B(n12473), .C(n11664), .D(n11325), 
        .Z(n8501) );
  HS65_LL_NAND2X2 U10987 ( .A(n10107), .B(n11746), .Z(n12506) );
  HS65_LL_NAND4ABX3 U10988 ( .A(n12469), .B(n12535), .C(n8501), .D(n12506), 
        .Z(n8509) );
  HS65_LL_IVX2 U10989 ( .A(sa22[2]), .Z(n8505) );
  HS65_LL_NOR2X2 U10990 ( .A(sa22[4]), .B(n8505), .Z(n12951) );
  HS65_LL_IVX2 U10991 ( .A(n8510), .Z(n8507) );
  HS65_LL_NAND2X2 U10992 ( .A(n10121), .B(n12501), .Z(n11764) );
  HS65_LL_NAND2X2 U10993 ( .A(n10123), .B(n12473), .Z(n12488) );
  HS65_LL_NAND2X2 U10994 ( .A(n8502), .B(n12929), .Z(n11313) );
  HS65_LL_NAND2X2 U10995 ( .A(n11322), .B(n11313), .Z(n12514) );
  HS65_LL_NAND4ABX3 U10996 ( .A(n12469), .B(n12514), .C(n12527), .D(n12449), 
        .Z(n8503) );
  HS65_LL_NOR3X1 U10997 ( .A(n11764), .B(n12488), .C(n8503), .Z(n12949) );
  HS65_LL_NOR2X2 U10998 ( .A(n12913), .B(n10127), .Z(n12459) );
  HS65_LL_IVX2 U10999 ( .A(n11323), .Z(n11311) );
  HS65_LL_NAND2X2 U11000 ( .A(n11311), .B(n10107), .Z(n11739) );
  HS65_LL_AND2X4 U11001 ( .A(n10116), .B(n11739), .Z(n12528) );
  HS65_LL_NOR4ABX2 U11002 ( .A(n12459), .B(n12528), .C(n12462), .D(n8504), .Z(
        n8506) );
  HS65_LL_NAND2X2 U11003 ( .A(sa22[4]), .B(n8505), .Z(n12947) );
  HS65_LL_AOI13X2 U11004 ( .A(n8507), .B(n12949), .C(n8506), .D(n12947), .Z(
        n8508) );
  HS65_LL_CBI4I6X2 U11005 ( .A(n8510), .B(n8509), .C(n12951), .D(n8508), .Z(
        n8511) );
  HS65_LL_CBI4I1X3 U11006 ( .A(n12495), .B(n8512), .C(n11339), .D(n8511), .Z(
        n8513) );
  HS65_LL_AOI12X2 U11007 ( .A(n12945), .B(n8514), .C(n8513), .Z(n15354) );
  HS65_LL_IVX2 U11008 ( .A(n15354), .Z(n15353) );
  HS65_LL_NOR2X2 U11009 ( .A(n13578), .B(n11207), .Z(n13960) );
  HS65_LL_NOR2X2 U11010 ( .A(n11200), .B(n13960), .Z(n11620) );
  HS65_LL_AOI112X2 U11011 ( .A(n8515), .B(n12976), .C(n13599), .D(n13598), .Z(
        n8523) );
  HS65_LL_NOR2X2 U11012 ( .A(n11208), .B(n11207), .Z(n12409) );
  HS65_LL_NAND2X2 U11013 ( .A(n8524), .B(n11635), .Z(n8519) );
  HS65_LL_NOR2X2 U11014 ( .A(n8516), .B(n12975), .Z(n13953) );
  HS65_LL_NOR4ABX2 U11015 ( .A(n12954), .B(n13953), .C(n8530), .D(n12997), .Z(
        n8518) );
  HS65_LL_NAND4ABX3 U11016 ( .A(n12409), .B(n8519), .C(n8518), .D(n8517), .Z(
        n12421) );
  HS65_LL_NOR2X2 U11017 ( .A(n8521), .B(n8520), .Z(n11641) );
  HS65_LL_NAND4ABX3 U11018 ( .A(n12960), .B(n11641), .C(n11630), .D(n13943), 
        .Z(n8522) );
  HS65_LL_NOR4ABX2 U11019 ( .A(n11620), .B(n8523), .C(n12421), .D(n8522), .Z(
        n8550) );
  HS65_LL_IVX2 U11020 ( .A(n13961), .Z(n12434) );
  HS65_LL_AND2X4 U11021 ( .A(n13585), .B(n13968), .Z(n11638) );
  HS65_LL_NOR4ABX2 U11022 ( .A(n8524), .B(n13593), .C(n12398), .D(n13960), .Z(
        n8525) );
  HS65_LL_NAND3X2 U11023 ( .A(n8526), .B(n11638), .C(n8525), .Z(n12969) );
  HS65_LL_IVX2 U11024 ( .A(n12996), .Z(n11204) );
  HS65_LL_NOR2X2 U11025 ( .A(n13602), .B(n11211), .Z(n12411) );
  HS65_LL_NOR2X2 U11026 ( .A(n11208), .B(n11623), .Z(n13574) );
  HS65_LL_NOR2X2 U11027 ( .A(n11641), .B(n13574), .Z(n11214) );
  HS65_LL_NAND2X2 U11028 ( .A(n11630), .B(n11646), .Z(n12998) );
  HS65_LL_NOR4ABX2 U11029 ( .A(n11214), .B(n12403), .C(n8527), .D(n12998), .Z(
        n8528) );
  HS65_LL_NAND4ABX3 U11030 ( .A(n12417), .B(n13575), .C(n12411), .D(n8528), 
        .Z(n13597) );
  HS65_LL_NAND2X2 U11031 ( .A(n8541), .B(n11203), .Z(n12407) );
  HS65_LL_NOR4ABX2 U11032 ( .A(n8536), .B(n11204), .C(n13597), .D(n12407), .Z(
        n8546) );
  HS65_LL_IVX2 U11033 ( .A(n13965), .Z(n12415) );
  HS65_LL_NOR4ABX2 U11034 ( .A(n12423), .B(n11635), .C(n12415), .D(n12962), 
        .Z(n8529) );
  HS65_LL_NAND4ABX3 U11035 ( .A(n11656), .B(n8530), .C(n8546), .D(n8529), .Z(
        n8548) );
  HS65_LL_NOR3X1 U11036 ( .A(n12416), .B(n12981), .C(n13966), .Z(n13573) );
  HS65_LL_NOR4ABX2 U11037 ( .A(n11195), .B(n13593), .C(n13599), .D(n13583), 
        .Z(n8532) );
  HS65_LL_NOR4ABX2 U11038 ( .A(n8532), .B(n8531), .C(n11644), .D(n13604), .Z(
        n11212) );
  HS65_LL_NAND3X2 U11039 ( .A(n8533), .B(n13943), .C(n12423), .Z(n8534) );
  HS65_LL_NOR4ABX2 U11040 ( .A(n12406), .B(n13585), .C(n12999), .D(n8534), .Z(
        n13964) );
  HS65_LL_NAND4ABX3 U11041 ( .A(n13576), .B(n12398), .C(n11212), .D(n13964), 
        .Z(n8535) );
  HS65_LL_NOR4ABX2 U11042 ( .A(n13573), .B(n12955), .C(n12409), .D(n8535), .Z(
        n8545) );
  HS65_LL_IVX2 U11043 ( .A(n13614), .Z(n13978) );
  HS65_LL_NAND2X2 U11044 ( .A(n8536), .B(n11201), .Z(n12978) );
  HS65_LL_NOR3X1 U11045 ( .A(n12412), .B(n12962), .C(n12998), .Z(n13582) );
  HS65_LL_IVX2 U11046 ( .A(n11202), .Z(n13603) );
  HS65_LL_NAND4ABX3 U11047 ( .A(n12960), .B(n13603), .C(n8537), .D(n12418), 
        .Z(n8538) );
  HS65_LL_NOR2X2 U11048 ( .A(n12990), .B(n12415), .Z(n11631) );
  HS65_LL_NAND4ABX3 U11049 ( .A(n13602), .B(n8538), .C(n11631), .D(n12410), 
        .Z(n13955) );
  HS65_LL_AOI112X2 U11050 ( .A(n11220), .B(n8539), .C(n12996), .D(n13955), .Z(
        n8540) );
  HS65_LL_NAND3X2 U11051 ( .A(n13573), .B(n8540), .C(n12403), .Z(n11196) );
  HS65_LL_NOR4ABX2 U11052 ( .A(n8541), .B(n11635), .C(n12417), .D(n11196), .Z(
        n8542) );
  HS65_LL_NAND4ABX3 U11053 ( .A(n13967), .B(n13568), .C(n13582), .D(n8542), 
        .Z(n8543) );
  HS65_LL_OAI13X1 U11054 ( .A(n13599), .B(n12978), .C(n8543), .D(n13981), .Z(
        n8544) );
  HS65_LL_CBI4I1X3 U11055 ( .A(n8546), .B(n8545), .C(n13978), .D(n8544), .Z(
        n8547) );
  HS65_LL_CBI4I6X2 U11056 ( .A(n12969), .B(n8548), .C(n13972), .D(n8547), .Z(
        n8549) );
  HS65_LL_CBI4I1X3 U11057 ( .A(n8551), .B(n8550), .C(n12434), .D(n8549), .Z(
        n15258) );
  HS65_LL_MUXI21X2 U11058 ( .D0(n15353), .D1(n15354), .S0(n15258), .Z(n14140)
         );
  HS65_LLS_XOR3X2 U11059 ( .A(n14819), .B(w0[26]), .C(n14140), .Z(n8552) );
  HS65_LLS_XOR3X2 U11060 ( .A(n15259), .B(n15552), .C(n8552), .Z(n8553) );
  HS65_LL_MUX31X4 U11061 ( .D0(w0[26]), .D1(n15120), .D2(n8553), .S0(
        text_in_r[122]), .S1(n14808), .Z(N276) );
  HS65_LL_IVX2 U11062 ( .A(w2[3]), .Z(n15509) );
  HS65_LL_NOR2AX3 U11063 ( .A(n8931), .B(n8940), .Z(n8729) );
  HS65_LL_NAND2X2 U11064 ( .A(n8554), .B(n8564), .Z(n15457) );
  HS65_LL_IVX2 U11065 ( .A(n15457), .Z(n8588) );
  HS65_LL_AOI12X2 U11066 ( .A(n8740), .B(n8739), .C(n8588), .Z(n15464) );
  HS65_LL_IVX2 U11067 ( .A(n12378), .Z(n12352) );
  HS65_LL_NAND3X2 U11068 ( .A(n15464), .B(n12352), .C(n8555), .Z(n8758) );
  HS65_LL_NAND2X2 U11069 ( .A(n8739), .B(n8563), .Z(n12351) );
  HS65_LL_NAND3X2 U11070 ( .A(n12371), .B(n12379), .C(n12351), .Z(n8556) );
  HS65_LL_NOR4ABX2 U11071 ( .A(n8557), .B(n8729), .C(n8758), .D(n8556), .Z(
        n13314) );
  HS65_LL_NOR2X2 U11072 ( .A(n8558), .B(n8902), .Z(n12377) );
  HS65_LL_NOR2X2 U11073 ( .A(n15485), .B(n12377), .Z(n8579) );
  HS65_LL_NAND3X2 U11074 ( .A(n8559), .B(n13314), .C(n8579), .Z(n8568) );
  HS65_LL_NOR2AX3 U11075 ( .A(n12363), .B(n12350), .Z(n8580) );
  HS65_LL_NAND2X2 U11076 ( .A(n8580), .B(n8560), .Z(n13331) );
  HS65_LL_NOR2X2 U11077 ( .A(n8561), .B(n8753), .Z(n8938) );
  HS65_LL_NAND4ABX3 U11078 ( .A(n15472), .B(n13331), .C(n8562), .D(n8938), .Z(
        n8760) );
  HS65_LL_NAND2X2 U11079 ( .A(n8909), .B(n8563), .Z(n15475) );
  HS65_LL_NAND3X2 U11080 ( .A(sa31[5]), .B(sa31[0]), .C(n13303), .Z(n13325) );
  HS65_LL_NAND3X2 U11081 ( .A(n15475), .B(n13325), .C(n13336), .Z(n15459) );
  HS65_LL_NOR2X2 U11082 ( .A(n8934), .B(n15459), .Z(n8925) );
  HS65_LL_NAND3X2 U11083 ( .A(sa31[1]), .B(n8564), .C(n12370), .Z(n13319) );
  HS65_LL_NAND2X2 U11084 ( .A(n15486), .B(n8749), .Z(n8900) );
  HS65_LL_NOR3X1 U11085 ( .A(n15489), .B(n13066), .C(n8900), .Z(n8566) );
  HS65_LL_NAND3X2 U11086 ( .A(n13319), .B(n8566), .C(n8565), .Z(n13080) );
  HS65_LL_NOR4ABX2 U11087 ( .A(n8723), .B(n8734), .C(n13311), .D(n13080), .Z(
        n8567) );
  HS65_LL_NAND4ABX3 U11088 ( .A(n8568), .B(n8760), .C(n8925), .D(n8567), .Z(
        n8595) );
  HS65_LL_IVX2 U11089 ( .A(n8568), .Z(n8576) );
  HS65_LL_NOR2X2 U11090 ( .A(n8569), .B(n12369), .Z(n8897) );
  HS65_LL_NAND3X2 U11091 ( .A(sa31[3]), .B(n8570), .C(n8739), .Z(n13317) );
  HS65_LL_NAND2X2 U11092 ( .A(n13317), .B(n8571), .Z(n12374) );
  HS65_LL_NOR3X1 U11093 ( .A(n12380), .B(n8897), .C(n12374), .Z(n8573) );
  HS65_LL_NAND2X2 U11094 ( .A(n8572), .B(n15482), .Z(n8922) );
  HS65_LL_NOR4ABX2 U11095 ( .A(n8573), .B(n13076), .C(n15489), .D(n8922), .Z(
        n8575) );
  HS65_LL_AOI13X2 U11096 ( .A(n8576), .B(n15460), .C(n8575), .D(n8574), .Z(
        n8594) );
  HS65_LL_NOR2X2 U11097 ( .A(n8930), .B(n13066), .Z(n8732) );
  HS65_LL_NAND3AX3 U11098 ( .A(n15459), .B(n13059), .C(n8732), .Z(n8577) );
  HS65_LL_NOR3X1 U11099 ( .A(n13305), .B(n8920), .C(n8577), .Z(n8748) );
  HS65_LL_NOR2X2 U11100 ( .A(n8897), .B(n8578), .Z(n8927) );
  HS65_LL_NOR2X2 U11101 ( .A(n15489), .B(n8737), .Z(n8757) );
  HS65_LL_NAND2X2 U11102 ( .A(n15464), .B(n8757), .Z(n13350) );
  HS65_LL_NAND4ABX3 U11103 ( .A(n13064), .B(n13350), .C(n8580), .D(n8579), .Z(
        n8581) );
  HS65_LL_NOR4ABX2 U11104 ( .A(n8927), .B(n13318), .C(n8932), .D(n8581), .Z(
        n8592) );
  HS65_LL_NOR4ABX2 U11105 ( .A(n8757), .B(n8583), .C(n12372), .D(n8582), .Z(
        n8584) );
  HS65_LL_NAND3X2 U11106 ( .A(n8584), .B(n8724), .C(n8749), .Z(n15505) );
  HS65_LL_NAND2X2 U11107 ( .A(n12381), .B(n15483), .Z(n8727) );
  HS65_LL_NOR2X2 U11108 ( .A(n8940), .B(n15484), .Z(n8923) );
  HS65_LL_IVX2 U11109 ( .A(n13303), .Z(n8756) );
  HS65_LL_NOR2X2 U11110 ( .A(n8585), .B(n8756), .Z(n8747) );
  HS65_LL_NAND2X2 U11111 ( .A(n13337), .B(n12363), .Z(n13056) );
  HS65_LL_NOR3X1 U11112 ( .A(n8747), .B(n13056), .C(n8586), .Z(n8587) );
  HS65_LL_NAND4ABX3 U11113 ( .A(n8588), .B(n8727), .C(n8923), .D(n8587), .Z(
        n8589) );
  HS65_LL_OAI13X1 U11114 ( .A(n8590), .B(n15505), .C(n8589), .D(n15494), .Z(
        n8591) );
  HS65_LL_CBI4I1X3 U11115 ( .A(n8748), .B(n8592), .C(n15500), .D(n8591), .Z(
        n8593) );
  HS65_LL_AOI112X2 U11116 ( .A(n15478), .B(n8595), .C(n8594), .D(n8593), .Z(
        n15510) );
  HS65_LL_NOR3AX2 U11117 ( .A(n8704), .B(n15171), .C(n8950), .Z(n8607) );
  HS65_LL_NAND4ABX3 U11118 ( .A(n9084), .B(n8596), .C(n8607), .D(n8613), .Z(
        n14483) );
  HS65_LL_NOR2X2 U11119 ( .A(n14475), .B(n8691), .Z(n9108) );
  HS65_LL_NOR4ABX2 U11120 ( .A(n9108), .B(n9089), .C(n8864), .D(n9118), .Z(
        n8597) );
  HS65_LL_NAND3X2 U11121 ( .A(n8717), .B(n8597), .C(n8684), .Z(n8679) );
  HS65_LL_NAND2AX4 U11122 ( .A(n8599), .B(n8598), .Z(n15144) );
  HS65_LL_NAND2X2 U11123 ( .A(n8956), .B(n8712), .Z(n8962) );
  HS65_LL_NAND2X2 U11124 ( .A(n15144), .B(n8962), .Z(n15167) );
  HS65_LL_NOR4ABX2 U11125 ( .A(n8951), .B(n8862), .C(n8877), .D(n9131), .Z(
        n8600) );
  HS65_LL_NAND3X2 U11126 ( .A(n8602), .B(n8601), .C(n8600), .Z(n8603) );
  HS65_LL_NOR3X1 U11127 ( .A(n8688), .B(n15167), .C(n8603), .Z(n9107) );
  HS65_LL_NOR2X2 U11128 ( .A(n14478), .B(n8972), .Z(n8614) );
  HS65_LL_NOR4ABX2 U11129 ( .A(n9107), .B(n8614), .C(n9092), .D(n8611), .Z(
        n8609) );
  HS65_LL_NOR2X2 U11130 ( .A(n8673), .B(n8695), .Z(n15159) );
  HS65_LL_NOR2X2 U11131 ( .A(n8673), .B(n8953), .Z(n9119) );
  HS65_LL_NOR3X1 U11132 ( .A(n8686), .B(n15159), .C(n9119), .Z(n15145) );
  HS65_LL_IVX2 U11133 ( .A(n8696), .Z(n8867) );
  HS65_LL_NOR3X1 U11134 ( .A(sa02[3]), .B(sa02[5]), .C(n8604), .Z(n15170) );
  HS65_LL_NOR4ABX2 U11135 ( .A(n15145), .B(n8867), .C(n8605), .D(n15170), .Z(
        n8606) );
  HS65_LL_NAND4ABX3 U11136 ( .A(n14483), .B(n8679), .C(n8609), .D(n8606), .Z(
        n8628) );
  HS65_LL_NOR2X2 U11137 ( .A(n9097), .B(n8871), .Z(n8850) );
  HS65_LL_NAND2X2 U11138 ( .A(n8852), .B(n9116), .Z(n14469) );
  HS65_LL_NOR4ABX2 U11139 ( .A(n8850), .B(n8607), .C(n8855), .D(n14469), .Z(
        n8608) );
  HS65_LL_NAND3X2 U11140 ( .A(n15147), .B(n8609), .C(n8608), .Z(n8627) );
  HS65_LL_OR3X4 U11141 ( .A(n15167), .B(n15171), .C(n8698), .Z(n9091) );
  HS65_LL_NOR2X2 U11142 ( .A(n8851), .B(n9091), .Z(n8682) );
  HS65_LL_NAND3X2 U11143 ( .A(n15145), .B(n14482), .C(n8862), .Z(n8610) );
  HS65_LL_AOI112X2 U11144 ( .A(n8958), .B(n8612), .C(n8611), .D(n8610), .Z(
        n8715) );
  HS65_LL_NAND2X2 U11145 ( .A(n9116), .B(n15154), .Z(n8866) );
  HS65_LL_NAND2X2 U11146 ( .A(n8613), .B(n15172), .Z(n9135) );
  HS65_LL_NOR4ABX2 U11147 ( .A(n8614), .B(n9108), .C(n8866), .D(n9135), .Z(
        n8615) );
  HS65_LL_NAND3X2 U11148 ( .A(n8682), .B(n8715), .C(n8615), .Z(n8626) );
  HS65_LL_NOR2X2 U11149 ( .A(n15171), .B(n8698), .Z(n8618) );
  HS65_LL_OR3X4 U11150 ( .A(n9125), .B(n8616), .C(n14478), .Z(n15175) );
  HS65_LL_NOR4ABX2 U11151 ( .A(n8618), .B(n8708), .C(n8617), .D(n15175), .Z(
        n15148) );
  HS65_LL_OAI21X2 U11152 ( .A(n8673), .B(n8619), .C(n8862), .Z(n8705) );
  HS65_LL_NOR3X1 U11153 ( .A(n14488), .B(n15149), .C(n8705), .Z(n8620) );
  HS65_LL_OAI112X1 U11154 ( .A(n8622), .B(n8621), .C(n15148), .D(n8620), .Z(
        n8623) );
  HS65_LL_IVX2 U11155 ( .A(n9123), .Z(n9096) );
  HS65_LL_NOR2X2 U11156 ( .A(n14475), .B(n9096), .Z(n9085) );
  HS65_LL_NOR2X2 U11157 ( .A(n8864), .B(n9100), .Z(n8954) );
  HS65_LL_NAND4ABX3 U11158 ( .A(n8624), .B(n8623), .C(n9085), .D(n8954), .Z(
        n8625) );
  HS65_LL_MX41X4 U11159 ( .D0(n8628), .S0(n15184), .D1(n8627), .S1(n15186), 
        .D2(n8626), .S2(n15182), .D3(n8625), .S3(n15180), .Z(n15629) );
  HS65_LLS_XNOR2X3 U11160 ( .A(n15510), .B(n15629), .Z(n15609) );
  HS65_LL_NAND2X2 U11161 ( .A(n8809), .B(n8630), .Z(n8662) );
  HS65_LL_NOR4ABX2 U11162 ( .A(n8837), .B(n8662), .C(n8841), .D(n12248), .Z(
        n8648) );
  HS65_LL_IVX2 U11163 ( .A(n8652), .Z(n15303) );
  HS65_LL_NAND2X2 U11164 ( .A(n8630), .B(n8629), .Z(n9018) );
  HS65_LL_NAND3X2 U11165 ( .A(n9018), .B(n12239), .C(n8805), .Z(n12262) );
  HS65_LL_NAND3X2 U11166 ( .A(n8657), .B(n8632), .C(n8631), .Z(n8633) );
  HS65_LL_NOR4X4 U11167 ( .A(n15303), .B(n12262), .C(n8634), .D(n8633), .Z(
        n8820) );
  HS65_LL_IVX2 U11168 ( .A(n8641), .Z(n8833) );
  HS65_LL_IVX2 U11169 ( .A(n12278), .Z(n12251) );
  HS65_LL_NAND3X2 U11170 ( .A(n8833), .B(n8992), .C(n12251), .Z(n15316) );
  HS65_LL_AOI12X2 U11171 ( .A(n8663), .B(n12264), .C(n15316), .Z(n8637) );
  HS65_LL_NAND2X2 U11172 ( .A(n8636), .B(n8635), .Z(n14502) );
  HS65_LL_NOR4ABX2 U11173 ( .A(n8820), .B(n8637), .C(n12247), .D(n14502), .Z(
        n8638) );
  HS65_LL_NAND3X2 U11174 ( .A(n8639), .B(n8648), .C(n8638), .Z(n8672) );
  HS65_LL_NAND4ABX3 U11175 ( .A(n8641), .B(n14515), .C(n8640), .D(n15305), .Z(
        n15292) );
  HS65_LL_NOR2X2 U11176 ( .A(n9002), .B(n8988), .Z(n8642) );
  HS65_LL_NOR3X1 U11177 ( .A(n12285), .B(n8643), .C(n8642), .Z(n8644) );
  HS65_LL_OAI21X2 U11178 ( .A(n15282), .B(n12274), .C(n8644), .Z(n8650) );
  HS65_LL_NOR2X2 U11179 ( .A(n14526), .B(n12244), .Z(n8666) );
  HS65_LL_NAND2X2 U11180 ( .A(n8645), .B(n8992), .Z(n15313) );
  HS65_LL_NOR3X1 U11181 ( .A(n8807), .B(n15313), .C(n8646), .Z(n8647) );
  HS65_LL_NAND3X2 U11182 ( .A(n8666), .B(n8648), .C(n8647), .Z(n14527) );
  HS65_LL_NOR2X2 U11183 ( .A(n8838), .B(n14527), .Z(n8826) );
  HS65_LL_NAND4ABX3 U11184 ( .A(n15292), .B(n8650), .C(n8826), .D(n8649), .Z(
        n8671) );
  HS65_LL_NAND3X2 U11185 ( .A(n9018), .B(n8651), .C(n12280), .Z(n12243) );
  HS65_LL_NAND4ABX3 U11186 ( .A(n12248), .B(n12243), .C(n8652), .D(n12239), 
        .Z(n8985) );
  HS65_LL_NOR2X2 U11187 ( .A(n8839), .B(n8653), .Z(n14501) );
  HS65_LL_OAI21X2 U11188 ( .A(n8988), .B(n9002), .C(n15299), .Z(n9027) );
  HS65_LL_NOR3X1 U11189 ( .A(n8655), .B(n8654), .C(n14506), .Z(n8656) );
  HS65_LL_NOR4ABX2 U11190 ( .A(n12271), .B(n8656), .C(n8807), .D(n15316), .Z(
        n14511) );
  HS65_LL_NAND4ABX3 U11191 ( .A(n8840), .B(n9027), .C(n8657), .D(n14511), .Z(
        n9017) );
  HS65_LL_NOR4ABX2 U11192 ( .A(n14501), .B(n15305), .C(n8658), .D(n9017), .Z(
        n8660) );
  HS65_LL_NAND4ABX3 U11193 ( .A(n8661), .B(n8985), .C(n8660), .D(n8659), .Z(
        n8670) );
  HS65_LL_NAND2X2 U11194 ( .A(n8842), .B(n8662), .Z(n9013) );
  HS65_LL_CBI4I6X2 U11195 ( .A(sa13[5]), .B(n8664), .C(n8663), .D(n9013), .Z(
        n8668) );
  HS65_LL_NOR4ABX2 U11196 ( .A(n8666), .B(n15315), .C(n14513), .D(n8665), .Z(
        n8667) );
  HS65_LL_NAND3X2 U11197 ( .A(n8668), .B(n8667), .C(n8822), .Z(n8669) );
  HS65_LL_MX41X4 U11198 ( .D0(n8672), .S0(n15328), .D1(n8671), .S1(n15326), 
        .D2(n8670), .S2(n15324), .D3(n8669), .S3(n15322), .Z(n15331) );
  HS65_LLS_XNOR2X3 U11199 ( .A(n15421), .B(n15331), .Z(n14627) );
  HS65_LL_NOR3X1 U11200 ( .A(n8675), .B(n8674), .C(n8673), .Z(n9105) );
  HS65_LL_NAND2X2 U11201 ( .A(n9111), .B(n8709), .Z(n15162) );
  HS65_LL_NAND3X2 U11202 ( .A(n15141), .B(n15162), .C(n8676), .Z(n8677) );
  HS65_LL_NOR3X1 U11203 ( .A(n9105), .B(n8678), .C(n8677), .Z(n15176) );
  HS65_LL_NOR4ABX2 U11204 ( .A(n8680), .B(n8951), .C(n9096), .D(n8679), .Z(
        n8681) );
  HS65_LL_NAND3X2 U11205 ( .A(n8682), .B(n15176), .C(n8681), .Z(n8722) );
  HS65_LL_NOR2AX3 U11206 ( .A(n8684), .B(n8683), .Z(n8861) );
  HS65_LL_NAND2AX4 U11207 ( .A(n9100), .B(n9101), .Z(n8685) );
  HS65_LL_NOR4ABX2 U11208 ( .A(n8687), .B(n8861), .C(n8686), .D(n8685), .Z(
        n8969) );
  HS65_LL_NOR3X1 U11209 ( .A(n15149), .B(n9124), .C(n8688), .Z(n8860) );
  HS65_LL_NAND4ABX3 U11210 ( .A(n15159), .B(n9098), .C(n8689), .D(n15162), .Z(
        n8690) );
  HS65_LL_NAND4ABX3 U11211 ( .A(n8866), .B(n8690), .C(n9083), .D(n9082), .Z(
        n8965) );
  HS65_LL_NOR4ABX2 U11212 ( .A(n8860), .B(n8692), .C(n8691), .D(n8965), .Z(
        n8693) );
  HS65_LL_NAND4ABX3 U11213 ( .A(n9091), .B(n14487), .C(n8969), .D(n8693), .Z(
        n8721) );
  HS65_LL_NOR2X2 U11214 ( .A(n8695), .B(n8694), .Z(n8876) );
  HS65_LL_NAND2X2 U11215 ( .A(n9122), .B(n9129), .Z(n8697) );
  HS65_LL_NOR2X2 U11216 ( .A(n8696), .B(n9120), .Z(n8849) );
  HS65_LL_NAND4ABX3 U11217 ( .A(n8876), .B(n8697), .C(n8849), .D(n8962), .Z(
        n14474) );
  HS65_LL_NOR3X1 U11218 ( .A(n8698), .B(n8950), .C(n15153), .Z(n8699) );
  HS65_LL_NAND3X2 U11219 ( .A(n8701), .B(n8700), .C(n8699), .Z(n8870) );
  HS65_LL_NOR2X2 U11220 ( .A(n15171), .B(n15149), .Z(n8703) );
  HS65_LL_NAND4ABX3 U11221 ( .A(n8859), .B(n8870), .C(n8703), .D(n8702), .Z(
        n8707) );
  HS65_LL_NOR2X2 U11222 ( .A(n8851), .B(n9098), .Z(n15173) );
  HS65_LL_NAND2X2 U11223 ( .A(n15173), .B(n8704), .Z(n14495) );
  HS65_LL_NOR4ABX2 U11224 ( .A(n8850), .B(n15144), .C(n8705), .D(n14495), .Z(
        n9114) );
  HS65_LL_NAND4ABX3 U11225 ( .A(n14474), .B(n8707), .C(n9114), .D(n8706), .Z(
        n8720) );
  HS65_LL_IVX2 U11226 ( .A(n8708), .Z(n8878) );
  HS65_LL_AOI12X2 U11227 ( .A(n8710), .B(n8709), .C(n8878), .Z(n8869) );
  HS65_LL_OAI21X2 U11228 ( .A(n8713), .B(n8712), .C(n8711), .Z(n9115) );
  HS65_LL_IVX2 U11229 ( .A(n8877), .Z(n8947) );
  HS65_LL_NAND2X2 U11230 ( .A(n8947), .B(n8714), .Z(n15160) );
  HS65_LL_IVX2 U11231 ( .A(n8876), .Z(n8966) );
  HS65_LL_NAND4ABX3 U11232 ( .A(n15161), .B(n15143), .C(n8715), .D(n8966), .Z(
        n8716) );
  HS65_LL_NOR4ABX2 U11233 ( .A(n8717), .B(n9115), .C(n15160), .D(n8716), .Z(
        n8718) );
  HS65_LL_NAND4ABX3 U11234 ( .A(n15171), .B(n9092), .C(n8869), .D(n8718), .Z(
        n8719) );
  HS65_LL_MX41X4 U11235 ( .D0(n8722), .S0(n15186), .D1(n8721), .S1(n15184), 
        .D2(n8720), .S2(n15182), .D3(n8719), .S3(n15180), .Z(n15594) );
  HS65_LL_IVX2 U11236 ( .A(n15594), .Z(n15593) );
  HS65_LL_IVX2 U11237 ( .A(n13304), .Z(n8731) );
  HS65_LL_NAND2X2 U11238 ( .A(n8723), .B(n8731), .Z(n13063) );
  HS65_LL_NAND4ABX3 U11239 ( .A(n13310), .B(n13063), .C(n8724), .D(n15475), 
        .Z(n8725) );
  HS65_LL_NAND4ABX3 U11240 ( .A(n13324), .B(n8725), .C(n8927), .D(n15469), .Z(
        n12384) );
  HS65_LL_NAND3X2 U11241 ( .A(n8938), .B(n12371), .C(n13306), .Z(n8726) );
  HS65_LL_NOR3AX2 U11242 ( .A(n13336), .B(n8727), .C(n8726), .Z(n12367) );
  HS65_LL_NOR4ABX2 U11243 ( .A(n13318), .B(n8729), .C(n8933), .D(n8728), .Z(
        n8730) );
  HS65_LL_NAND4ABX3 U11244 ( .A(n13350), .B(n8735), .C(n12367), .D(n8730), .Z(
        n8765) );
  HS65_LL_NOR2X2 U11245 ( .A(n8747), .B(n8922), .Z(n8914) );
  HS65_LL_NAND2X2 U11246 ( .A(n15457), .B(n8731), .Z(n13073) );
  HS65_LL_NOR4ABX2 U11247 ( .A(n8732), .B(n8914), .C(n13064), .D(n13073), .Z(
        n13327) );
  HS65_LL_NOR2X2 U11248 ( .A(n8733), .B(n8745), .Z(n15466) );
  HS65_LL_NAND4ABX3 U11249 ( .A(n15466), .B(n8735), .C(n12348), .D(n8734), .Z(
        n8736) );
  HS65_LL_NOR3X1 U11250 ( .A(n12380), .B(n8737), .C(n8736), .Z(n13334) );
  HS65_LL_NAND3X2 U11251 ( .A(n13318), .B(n13317), .C(n12381), .Z(n8928) );
  HS65_LL_NOR2X2 U11252 ( .A(n8738), .B(n12359), .Z(n12366) );
  HS65_LL_AOI12X2 U11253 ( .A(n8740), .B(n8739), .C(n12366), .Z(n12349) );
  HS65_LL_NAND4ABX3 U11254 ( .A(n15484), .B(n8928), .C(n12349), .D(n8741), .Z(
        n13057) );
  HS65_LL_NAND4ABX3 U11255 ( .A(n8929), .B(n13057), .C(n8743), .D(n8742), .Z(
        n8744) );
  HS65_LL_NOR4ABX2 U11256 ( .A(n13327), .B(n13334), .C(n8940), .D(n8744), .Z(
        n8763) );
  HS65_LL_AOI12X2 U11257 ( .A(n8746), .B(n8745), .C(n12376), .Z(n8752) );
  HS65_LL_IVX2 U11258 ( .A(n12371), .Z(n15465) );
  HS65_LL_NOR3X1 U11259 ( .A(n12362), .B(n15465), .C(n12366), .Z(n8898) );
  HS65_LL_NAND2AX4 U11260 ( .A(n15493), .B(n12351), .Z(n13329) );
  HS65_LL_NOR4ABX2 U11261 ( .A(n8748), .B(n8898), .C(n8747), .D(n13329), .Z(
        n8750) );
  HS65_LL_NAND4ABX3 U11262 ( .A(n15466), .B(n15462), .C(n8750), .D(n8749), .Z(
        n8751) );
  HS65_LL_OAI13X1 U11263 ( .A(n8753), .B(n8752), .C(n8751), .D(n15494), .Z(
        n8762) );
  HS65_LL_NOR4ABX2 U11264 ( .A(n8754), .B(n12379), .C(n8919), .D(n8929), .Z(
        n8755) );
  HS65_LL_OAI21X2 U11265 ( .A(n8907), .B(n8756), .C(n8755), .Z(n15496) );
  HS65_LL_OR3X4 U11266 ( .A(n8933), .B(n13067), .C(n12372), .Z(n13330) );
  HS65_LL_NAND4ABX3 U11267 ( .A(n8758), .B(n13330), .C(n8911), .D(n8757), .Z(
        n8759) );
  HS65_LL_OAI13X1 U11268 ( .A(n15496), .B(n8760), .C(n8759), .D(n15503), .Z(
        n8761) );
  HS65_LL_OAI112X1 U11269 ( .A(n8763), .B(n15500), .C(n8762), .D(n8761), .Z(
        n8764) );
  HS65_LL_CBI4I6X2 U11270 ( .A(n12384), .B(n8765), .C(n15478), .D(n8764), .Z(
        n15455) );
  HS65_LL_MUXI21X2 U11271 ( .D0(n15594), .D1(n15593), .S0(n15455), .Z(n15624)
         );
  HS65_LLS_XOR3X2 U11272 ( .A(w2[3]), .B(n15624), .C(n15189), .Z(n8766) );
  HS65_LLS_XOR3X2 U11273 ( .A(n15609), .B(n14627), .C(n8766), .Z(n8767) );
  HS65_LL_MUXI31X2 U11274 ( .D0(n15509), .D1(w2[3]), .D2(n8767), .S0(
        text_in_r[35]), .S1(n14808), .Z(N101) );
  HS65_LL_IVX2 U11275 ( .A(w2[1]), .Z(n15512) );
  HS65_LL_NOR4ABX2 U11276 ( .A(n8769), .B(n8794), .C(n12310), .D(n8768), .Z(
        n8770) );
  HS65_LL_NAND4ABX3 U11277 ( .A(n12308), .B(n8772), .C(n8771), .D(n8770), .Z(
        n8804) );
  HS65_LL_NAND4ABX3 U11278 ( .A(n8774), .B(n8773), .C(n15396), .D(n13023), .Z(
        n13042) );
  HS65_LL_NAND3AX3 U11279 ( .A(n8776), .B(n8775), .C(n13032), .Z(n8777) );
  HS65_LL_NOR3X1 U11280 ( .A(n8779), .B(n8778), .C(n8777), .Z(n12328) );
  HS65_LL_NOR2X2 U11281 ( .A(n8800), .B(n8780), .Z(n15378) );
  HS65_LL_NAND2X2 U11282 ( .A(n15378), .B(n9047), .Z(n15399) );
  HS65_LL_NOR4ABX2 U11283 ( .A(n8782), .B(n12313), .C(n8781), .D(n15399), .Z(
        n8783) );
  HS65_LL_NAND4ABX3 U11284 ( .A(n8798), .B(n13042), .C(n12328), .D(n8783), .Z(
        n8803) );
  HS65_LL_NAND3X2 U11285 ( .A(sa20[6]), .B(n8785), .C(n8784), .Z(n12331) );
  HS65_LL_NAND2X2 U11286 ( .A(n9047), .B(n12331), .Z(n15375) );
  HS65_LL_NOR3X1 U11287 ( .A(n9071), .B(n12301), .C(n15375), .Z(n8790) );
  HS65_LL_NOR3X1 U11288 ( .A(n8787), .B(n8786), .C(n9065), .Z(n8789) );
  HS65_LL_NAND3X2 U11289 ( .A(n8789), .B(n13017), .C(n8788), .Z(n15402) );
  HS65_LL_NOR4ABX2 U11290 ( .A(n8790), .B(n15374), .C(n9033), .D(n15402), .Z(
        n8791) );
  HS65_LL_NAND3X2 U11291 ( .A(n9057), .B(n8792), .C(n8791), .Z(n8802) );
  HS65_LL_IVX2 U11292 ( .A(n8793), .Z(n13022) );
  HS65_LL_NOR2X2 U11293 ( .A(n13022), .B(n9075), .Z(n12326) );
  HS65_LL_NAND2X2 U11294 ( .A(n12326), .B(n8794), .Z(n15388) );
  HS65_LL_NAND3AX3 U11295 ( .A(n9044), .B(n8796), .C(n8795), .Z(n13050) );
  HS65_LL_NOR3X1 U11296 ( .A(n8798), .B(n13050), .C(n8797), .Z(n8799) );
  HS65_LL_NAND4ABX3 U11297 ( .A(n8800), .B(n15388), .C(n12337), .D(n8799), .Z(
        n8801) );
  HS65_LL_MX41X4 U11298 ( .D0(n8804), .S0(n13020), .D1(n8803), .S1(n15416), 
        .D2(n8802), .S2(n15408), .D3(n8801), .S3(n15400), .Z(n15425) );
  HS65_LL_NAND3X2 U11299 ( .A(n12237), .B(n8805), .C(n15299), .Z(n8806) );
  HS65_LL_NOR3AX2 U11300 ( .A(n15290), .B(n8807), .C(n8806), .Z(n15288) );
  HS65_LL_NOR2X2 U11301 ( .A(n12247), .B(n8838), .Z(n9019) );
  HS65_LL_NAND3X2 U11302 ( .A(sa13[6]), .B(n8809), .C(n8808), .Z(n15314) );
  HS65_LL_NAND2X2 U11303 ( .A(n8810), .B(n15314), .Z(n12238) );
  HS65_LL_NOR4ABX2 U11304 ( .A(n15288), .B(n9019), .C(n12283), .D(n12238), .Z(
        n8811) );
  HS65_LL_NAND4ABX3 U11305 ( .A(n8812), .B(n9005), .C(n15318), .D(n8811), .Z(
        n8848) );
  HS65_LL_NAND2X2 U11306 ( .A(n8813), .B(n15278), .Z(n14528) );
  HS65_LL_AOI12X2 U11307 ( .A(n8816), .B(n8815), .C(n8814), .Z(n15307) );
  HS65_LL_AOI12X2 U11308 ( .A(n8818), .B(n8817), .C(n15307), .Z(n8819) );
  HS65_LL_OAI21X2 U11309 ( .A(sa13[6]), .B(n12274), .C(n8819), .Z(n8821) );
  HS65_LL_NAND4ABX3 U11310 ( .A(n14528), .B(n8821), .C(n8828), .D(n8820), .Z(
        n8847) );
  HS65_LL_NAND2AX4 U11311 ( .A(n15280), .B(n8822), .Z(n14503) );
  HS65_LL_NOR2X2 U11312 ( .A(n14516), .B(n14503), .Z(n12286) );
  HS65_LL_NOR4ABX2 U11313 ( .A(n8824), .B(n12286), .C(n14514), .D(n8823), .Z(
        n8825) );
  HS65_LL_NAND3X2 U11314 ( .A(n8827), .B(n8826), .C(n8825), .Z(n8846) );
  HS65_LL_IVX2 U11315 ( .A(n8828), .Z(n8844) );
  HS65_LL_NOR2X2 U11316 ( .A(n9002), .B(n14522), .Z(n15285) );
  HS65_LL_NOR3X1 U11317 ( .A(n14533), .B(n15285), .C(n8829), .Z(n8830) );
  HS65_LL_OAI21X2 U11318 ( .A(n8990), .B(n8831), .C(n8830), .Z(n14519) );
  HS65_LL_NOR2X2 U11319 ( .A(n14522), .B(n8832), .Z(n8836) );
  HS65_LL_NAND3X2 U11320 ( .A(n8834), .B(n8833), .C(n9001), .Z(n8835) );
  HS65_LL_NOR3X1 U11321 ( .A(n8836), .B(n12259), .C(n8835), .Z(n12256) );
  HS65_LL_IVX2 U11322 ( .A(n8837), .Z(n14510) );
  HS65_LL_NOR3X1 U11323 ( .A(n14510), .B(n8839), .C(n8838), .Z(n15319) );
  HS65_LL_NAND2AX4 U11324 ( .A(n8840), .B(n9018), .Z(n12284) );
  HS65_LL_NOR4ABX2 U11325 ( .A(n15319), .B(n8842), .C(n8841), .D(n12284), .Z(
        n8843) );
  HS65_LL_NAND4ABX3 U11326 ( .A(n8844), .B(n14519), .C(n12256), .D(n8843), .Z(
        n8845) );
  HS65_LL_MX41X4 U11327 ( .D0(n8848), .S0(n15326), .D1(n8847), .S1(n15328), 
        .D2(n8846), .S2(n15324), .D3(n8845), .S3(n15322), .Z(n15334) );
  HS65_LLS_XOR2X3 U11328 ( .A(n15425), .B(n15334), .Z(n14946) );
  HS65_LL_NAND3X2 U11329 ( .A(n8850), .B(n15145), .C(n8849), .Z(n8896) );
  HS65_LL_NOR4ABX2 U11330 ( .A(n8853), .B(n8852), .C(n14477), .D(n8851), .Z(
        n8949) );
  HS65_LL_IVX2 U11331 ( .A(n9099), .Z(n14467) );
  HS65_LL_OR2X4 U11332 ( .A(n15149), .B(n9088), .Z(n8880) );
  HS65_LL_NAND4ABX3 U11333 ( .A(n8855), .B(n14488), .C(n8854), .D(n9083), .Z(
        n15152) );
  HS65_LL_NOR4ABX2 U11334 ( .A(n8949), .B(n14467), .C(n8880), .D(n15152), .Z(
        n8856) );
  HS65_LL_NAND4ABX3 U11335 ( .A(n9100), .B(n9118), .C(n8857), .D(n8856), .Z(
        n8895) );
  HS65_LL_NOR2X2 U11336 ( .A(n14475), .B(n8870), .Z(n9127) );
  HS65_LL_NAND2X2 U11337 ( .A(n9127), .B(n8858), .Z(n8974) );
  HS65_LL_NOR4ABX2 U11338 ( .A(n8861), .B(n8860), .C(n8859), .D(n8974), .Z(
        n8893) );
  HS65_LL_NAND2X2 U11339 ( .A(n8862), .B(n8868), .Z(n14468) );
  HS65_LL_NOR2X2 U11340 ( .A(n9121), .B(n8972), .Z(n8967) );
  HS65_LL_NOR4ABX2 U11341 ( .A(n9129), .B(n15144), .C(n8864), .D(n8863), .Z(
        n8865) );
  HS65_LL_NAND4ABX3 U11342 ( .A(n8971), .B(n8866), .C(n8967), .D(n8865), .Z(
        n15174) );
  HS65_LL_NOR4ABX2 U11343 ( .A(n8867), .B(n8966), .C(n14468), .D(n15174), .Z(
        n8892) );
  HS65_LL_NAND2AX4 U11344 ( .A(n9097), .B(n8868), .Z(n9086) );
  HS65_LL_NAND4ABX3 U11345 ( .A(n9096), .B(n9086), .C(n8869), .D(n15162), .Z(
        n8874) );
  HS65_LL_NAND4ABX3 U11346 ( .A(n9100), .B(n8870), .C(n14476), .D(n15145), .Z(
        n8873) );
  HS65_LL_NOR2X2 U11347 ( .A(n14488), .B(n8871), .Z(n8872) );
  HS65_LL_NAND4ABX3 U11348 ( .A(n8874), .B(n8873), .C(n9107), .D(n8872), .Z(
        n8889) );
  HS65_LL_NAND3X2 U11349 ( .A(sa02[6]), .B(n9111), .C(n8875), .Z(n15139) );
  HS65_LL_NOR3X1 U11350 ( .A(n8973), .B(n8877), .C(n8876), .Z(n9117) );
  HS65_LL_NAND4ABX3 U11351 ( .A(n8878), .B(n9121), .C(n15176), .D(n9117), .Z(
        n8879) );
  HS65_LL_NOR4ABX2 U11352 ( .A(n8881), .B(n15139), .C(n8880), .D(n8879), .Z(
        n14494) );
  HS65_LL_NOR3X1 U11353 ( .A(n9125), .B(n15159), .C(n8882), .Z(n8885) );
  HS65_LL_NAND2X2 U11354 ( .A(n8883), .B(n9082), .Z(n9104) );
  HS65_LL_NOR4ABX2 U11355 ( .A(n8885), .B(n8962), .C(n8884), .D(n9104), .Z(
        n8886) );
  HS65_LL_NAND3X2 U11356 ( .A(n8887), .B(n14494), .C(n8886), .Z(n8888) );
  HS65_LL_AOI22X1 U11357 ( .A(n15180), .B(n8889), .C(n15184), .D(n8888), .Z(
        n8890) );
  HS65_LL_CBI4I1X3 U11358 ( .A(n8893), .B(n8892), .C(n8891), .D(n8890), .Z(
        n8894) );
  HS65_LL_CBI4I6X2 U11359 ( .A(n8896), .B(n8895), .C(n15182), .D(n8894), .Z(
        n15625) );
  HS65_LL_NAND2AX4 U11360 ( .A(n13310), .B(n13317), .Z(n8905) );
  HS65_LL_IVX2 U11361 ( .A(n8897), .Z(n8918) );
  HS65_LL_NAND2X2 U11362 ( .A(n8898), .B(n8918), .Z(n13338) );
  HS65_LL_NOR2X2 U11363 ( .A(n13324), .B(n15458), .Z(n12365) );
  HS65_LL_NAND4ABX3 U11364 ( .A(n13305), .B(n8900), .C(n12365), .D(n8899), .Z(
        n8901) );
  HS65_LL_NOR3X1 U11365 ( .A(n15496), .B(n13338), .C(n8901), .Z(n13065) );
  HS65_LL_CBI4I1X3 U11366 ( .A(n8903), .B(n8902), .C(sa31[7]), .D(n13065), .Z(
        n8904) );
  HS65_LL_AOI112X2 U11367 ( .A(n8907), .B(n8906), .C(n8905), .D(n8904), .Z(
        n8908) );
  HS65_LL_NAND3X2 U11368 ( .A(n13348), .B(n8908), .C(n13347), .Z(n8944) );
  HS65_LL_NAND2X2 U11369 ( .A(n8910), .B(n8909), .Z(n12356) );
  HS65_LL_IVX2 U11370 ( .A(n15483), .Z(n13339) );
  HS65_LL_NAND4ABX3 U11371 ( .A(n13339), .B(n15459), .C(n13337), .D(n8911), 
        .Z(n8912) );
  HS65_LL_NOR4ABX2 U11372 ( .A(n8914), .B(n12356), .C(n8913), .D(n8912), .Z(
        n8915) );
  HS65_LL_NAND3X2 U11373 ( .A(n13314), .B(n13334), .C(n8915), .Z(n8943) );
  HS65_LL_NAND3X2 U11374 ( .A(n8917), .B(n13317), .C(n8916), .Z(n15481) );
  HS65_LL_NOR3X1 U11375 ( .A(n13305), .B(n12350), .C(n13310), .Z(n12358) );
  HS65_LL_NAND2X2 U11376 ( .A(n12358), .B(n8918), .Z(n13074) );
  HS65_LL_NOR3X1 U11377 ( .A(n8920), .B(n13064), .C(n8919), .Z(n8921) );
  HS65_LL_NAND3X2 U11378 ( .A(n8921), .B(n13076), .C(n15483), .Z(n12383) );
  HS65_LL_NOR4ABX2 U11379 ( .A(n8923), .B(n13344), .C(n8922), .D(n12383), .Z(
        n8924) );
  HS65_LL_NAND4ABX3 U11380 ( .A(n15481), .B(n13074), .C(n8925), .D(n8924), .Z(
        n8942) );
  HS65_LL_NOR4ABX2 U11381 ( .A(n12357), .B(n15457), .C(n12377), .D(n12347), 
        .Z(n8926) );
  HS65_LL_NAND4ABX3 U11382 ( .A(n13324), .B(n8928), .C(n8927), .D(n8926), .Z(
        n15497) );
  HS65_LL_NOR2X2 U11383 ( .A(n8930), .B(n8929), .Z(n8937) );
  HS65_LL_NAND4ABX3 U11384 ( .A(n8933), .B(n8932), .C(n8931), .D(n13347), .Z(
        n8936) );
  HS65_LL_NAND4ABX3 U11385 ( .A(n8934), .B(n12366), .C(n12363), .D(n15475), 
        .Z(n8935) );
  HS65_LL_NOR4ABX2 U11386 ( .A(n8938), .B(n8937), .C(n8936), .D(n8935), .Z(
        n8939) );
  HS65_LL_NAND4ABX3 U11387 ( .A(n8940), .B(n15497), .C(n13334), .D(n8939), .Z(
        n8941) );
  HS65_LL_MX41X4 U11388 ( .D0(n8944), .S0(n15478), .D1(n8943), .S1(n15494), 
        .D2(n8942), .S2(n13352), .D3(n8941), .S3(n15503), .Z(n15561) );
  HS65_LLS_XNOR2X3 U11389 ( .A(n15625), .B(n15561), .Z(n15600) );
  HS65_LL_NOR3X1 U11390 ( .A(n9125), .B(n9119), .C(n8945), .Z(n8948) );
  HS65_LL_NOR4ABX2 U11391 ( .A(n8948), .B(n8947), .C(n8973), .D(n8946), .Z(
        n14485) );
  HS65_LL_NAND4ABX3 U11392 ( .A(n8950), .B(n14468), .C(n8949), .D(n14485), .Z(
        n8955) );
  HS65_LL_OAI21X2 U11393 ( .A(n8953), .B(n8952), .C(n8951), .Z(n14473) );
  HS65_LL_NOR2X2 U11394 ( .A(n8972), .B(n14473), .Z(n15140) );
  HS65_LL_NAND4ABX3 U11395 ( .A(n8965), .B(n8955), .C(n8954), .D(n15140), .Z(
        n8980) );
  HS65_LL_NAND2X2 U11396 ( .A(sa02[1]), .B(n8956), .Z(n8960) );
  HS65_LL_NAND2X2 U11397 ( .A(n8958), .B(n8957), .Z(n8959) );
  HS65_LL_OAI112X1 U11398 ( .A(sa02[6]), .B(n8960), .C(n9115), .D(n8959), .Z(
        n8964) );
  HS65_LL_NOR4ABX2 U11399 ( .A(n8966), .B(n8962), .C(n8961), .D(n15153), .Z(
        n14471) );
  HS65_LL_NAND4ABX3 U11400 ( .A(n8965), .B(n8964), .C(n14471), .D(n8963), .Z(
        n8979) );
  HS65_LL_NAND3X2 U11401 ( .A(n8967), .B(n15139), .C(n8966), .Z(n8968) );
  HS65_LL_NOR4ABX2 U11402 ( .A(n8969), .B(n9082), .C(n15152), .D(n8968), .Z(
        n8970) );
  HS65_LL_NAND3X2 U11403 ( .A(n15148), .B(n9114), .C(n8970), .Z(n8978) );
  HS65_LL_NOR3X1 U11404 ( .A(n9099), .B(n8971), .C(n9118), .Z(n14489) );
  HS65_LL_NOR2X2 U11405 ( .A(n8973), .B(n8972), .Z(n15155) );
  HS65_LL_NOR4ABX2 U11406 ( .A(n15155), .B(n8975), .C(n9131), .D(n8974), .Z(
        n8976) );
  HS65_LL_NAND3X2 U11407 ( .A(n14466), .B(n14489), .C(n8976), .Z(n8977) );
  HS65_LL_MX41X4 U11408 ( .D0(n8980), .S0(n15186), .D1(n8979), .S1(n15184), 
        .D2(n8978), .S2(n15182), .D3(n8977), .S3(n15180), .Z(n15192) );
  HS65_LLS_XOR3X2 U11409 ( .A(n15624), .B(w2[1]), .C(n15192), .Z(n8981) );
  HS65_LLS_XOR3X2 U11410 ( .A(n14946), .B(n15600), .C(n8981), .Z(n8982) );
  HS65_LL_MUX31X4 U11411 ( .D0(w2[1]), .D1(n15512), .D2(n8982), .S0(
        text_in_r[33]), .S1(n14808), .Z(N99) );
  HS65_LL_IVX2 U11412 ( .A(w2[4]), .Z(n15507) );
  HS65_LL_NOR3X1 U11413 ( .A(n14526), .B(n12247), .C(n8983), .Z(n8984) );
  HS65_LL_NAND4ABX3 U11414 ( .A(n14514), .B(n8985), .C(n8984), .D(n12237), .Z(
        n8986) );
  HS65_LL_NOR3X1 U11415 ( .A(n12259), .B(n8987), .C(n8986), .Z(n15295) );
  HS65_LL_AOI112X2 U11416 ( .A(sa13[5]), .B(n8990), .C(n8989), .D(n8988), .Z(
        n8991) );
  HS65_LL_NOR4ABX2 U11417 ( .A(n8993), .B(n8992), .C(n8991), .D(n12265), .Z(
        n8994) );
  HS65_LL_NAND4ABX3 U11418 ( .A(n12257), .B(n14503), .C(n15295), .D(n8994), 
        .Z(n9031) );
  HS65_LL_NOR2X2 U11419 ( .A(n8996), .B(n8995), .Z(n8999) );
  HS65_LL_AOI112X2 U11420 ( .A(sa13[0]), .B(n8999), .C(n8998), .D(n8997), .Z(
        n9011) );
  HS65_LL_IVX2 U11421 ( .A(n9000), .Z(n9003) );
  HS65_LL_OAI21X2 U11422 ( .A(n9003), .B(n9002), .C(n9001), .Z(n9004) );
  HS65_LL_NOR3X1 U11423 ( .A(n15307), .B(n9005), .C(n9004), .Z(n15287) );
  HS65_LL_NOR4ABX2 U11424 ( .A(n9008), .B(n9007), .C(n12283), .D(n9006), .Z(
        n12242) );
  HS65_LL_NOR4ABX2 U11425 ( .A(n15287), .B(n12242), .C(n12288), .D(n9009), .Z(
        n9010) );
  HS65_LL_NAND3X2 U11426 ( .A(n12250), .B(n9011), .C(n9010), .Z(n9030) );
  HS65_LL_NAND4ABX3 U11427 ( .A(n9014), .B(n9013), .C(n12242), .D(n9012), .Z(
        n9016) );
  HS65_LL_NAND4ABX3 U11428 ( .A(n9017), .B(n9016), .C(n9015), .D(n12237), .Z(
        n9029) );
  HS65_LL_AND3X4 U11429 ( .A(n9020), .B(n9019), .C(n9018), .Z(n9021) );
  HS65_LL_NAND4ABX3 U11430 ( .A(n9022), .B(n15316), .C(n9021), .D(n12242), .Z(
        n9023) );
  HS65_LL_NOR4ABX2 U11431 ( .A(n9024), .B(n12260), .C(n12257), .D(n9023), .Z(
        n9026) );
  HS65_LL_NAND4ABX3 U11432 ( .A(n12240), .B(n9027), .C(n9026), .D(n9025), .Z(
        n9028) );
  HS65_LL_MX41X4 U11433 ( .D0(n9031), .S0(n15328), .D1(n9030), .S1(n15326), 
        .D2(n9029), .S2(n15324), .D3(n9028), .S3(n15322), .Z(n15569) );
  HS65_LL_NOR4ABX2 U11434 ( .A(n9035), .B(n9034), .C(n9033), .D(n9032), .Z(
        n12334) );
  HS65_LL_AOI12X2 U11435 ( .A(n9037), .B(n9036), .C(n13022), .Z(n9040) );
  HS65_LL_NOR4ABX2 U11436 ( .A(n9041), .B(n9040), .C(n9039), .D(n9038), .Z(
        n9042) );
  HS65_LL_NAND4ABX3 U11437 ( .A(n15376), .B(n9043), .C(n12334), .D(n9042), .Z(
        n9081) );
  HS65_LL_NOR4ABX2 U11438 ( .A(n12297), .B(n15381), .C(n9044), .D(n12323), .Z(
        n9052) );
  HS65_LL_NAND3X2 U11439 ( .A(n9046), .B(n9045), .C(n12313), .Z(n12335) );
  HS65_LL_NAND3X2 U11440 ( .A(n15377), .B(n13036), .C(n9047), .Z(n9048) );
  HS65_LL_NOR4ABX2 U11441 ( .A(n9049), .B(n12334), .C(n12335), .D(n9048), .Z(
        n9051) );
  HS65_LL_NAND3X2 U11442 ( .A(n9052), .B(n9051), .C(n9050), .Z(n9080) );
  HS65_LL_NOR3X1 U11443 ( .A(n9055), .B(n9054), .C(n9053), .Z(n9056) );
  HS65_LL_NAND3X2 U11444 ( .A(n9057), .B(n9056), .C(n13032), .Z(n15398) );
  HS65_LL_NAND3X2 U11445 ( .A(n9059), .B(n9058), .C(n12318), .Z(n9064) );
  HS65_LL_NOR4ABX2 U11446 ( .A(n9062), .B(n13023), .C(n9061), .D(n9060), .Z(
        n9063) );
  HS65_LL_NAND4ABX3 U11447 ( .A(n15398), .B(n9064), .C(n12334), .D(n9063), .Z(
        n9079) );
  HS65_LL_IVX2 U11448 ( .A(n9065), .Z(n12336) );
  HS65_LL_NAND2X2 U11449 ( .A(n9066), .B(n13016), .Z(n15383) );
  HS65_LL_NOR4ABX2 U11450 ( .A(n12336), .B(n9068), .C(n9067), .D(n15383), .Z(
        n9069) );
  HS65_LL_NAND4ABX3 U11451 ( .A(n9071), .B(n13034), .C(n9070), .D(n9069), .Z(
        n15406) );
  HS65_LL_NAND4ABX3 U11452 ( .A(n9073), .B(n12299), .C(n9072), .D(n15392), .Z(
        n9077) );
  HS65_LL_NOR3X1 U11453 ( .A(n12308), .B(n9075), .C(n9074), .Z(n13033) );
  HS65_LL_NAND4ABX3 U11454 ( .A(n15406), .B(n9077), .C(n9076), .D(n13033), .Z(
        n9078) );
  HS65_LL_MX41X4 U11455 ( .D0(n9081), .S0(n13020), .D1(n9080), .S1(n15416), 
        .D2(n9079), .S2(n15408), .D3(n9078), .S3(n15400), .Z(n15419) );
  HS65_LLS_XOR2X3 U11456 ( .A(n15569), .B(n15419), .Z(n15583) );
  HS65_LL_NAND2X2 U11457 ( .A(n9083), .B(n9082), .Z(n9087) );
  HS65_LL_NOR2X2 U11458 ( .A(n9100), .B(n9084), .Z(n15169) );
  HS65_LL_NAND4ABX3 U11459 ( .A(n9087), .B(n9086), .C(n9085), .D(n15169), .Z(
        n9095) );
  HS65_LL_NOR2X2 U11460 ( .A(n9088), .B(n15143), .Z(n9090) );
  HS65_LL_NAND4ABX3 U11461 ( .A(n9092), .B(n9091), .C(n9090), .D(n9089), .Z(
        n9094) );
  HS65_LL_NAND4ABX3 U11462 ( .A(n9095), .B(n9094), .C(n9093), .D(n9117), .Z(
        n9139) );
  HS65_LL_NOR3X1 U11463 ( .A(n9097), .B(n9096), .C(n15159), .Z(n14480) );
  HS65_LL_IVX2 U11464 ( .A(n9098), .Z(n14484) );
  HS65_LL_NOR4ABX2 U11465 ( .A(n9102), .B(n9101), .C(n9100), .D(n9099), .Z(
        n9103) );
  HS65_LL_NAND4ABX3 U11466 ( .A(n9105), .B(n9104), .C(n14484), .D(n9103), .Z(
        n15166) );
  HS65_LL_NOR4ABX2 U11467 ( .A(n9108), .B(n9107), .C(n9106), .D(n15166), .Z(
        n9109) );
  HS65_LL_NAND3X2 U11468 ( .A(n9110), .B(n14480), .C(n9109), .Z(n9138) );
  HS65_LL_AOI12X2 U11469 ( .A(n9112), .B(n9111), .C(n14477), .Z(n9113) );
  HS65_LL_NAND3X2 U11470 ( .A(n9115), .B(n9114), .C(n9113), .Z(n15158) );
  HS65_LL_NAND2X2 U11471 ( .A(n9117), .B(n9116), .Z(n9130) );
  HS65_LL_NOR2X2 U11472 ( .A(n9119), .B(n9118), .Z(n14470) );
  HS65_LL_NOR4ABX2 U11473 ( .A(n9123), .B(n9122), .C(n9121), .D(n9120), .Z(
        n9126) );
  HS65_LL_NOR4ABX2 U11474 ( .A(n9127), .B(n9126), .C(n9125), .D(n9124), .Z(
        n9128) );
  HS65_LL_NAND4ABX3 U11475 ( .A(n15158), .B(n9130), .C(n14470), .D(n9128), .Z(
        n9137) );
  HS65_LL_NAND4ABX3 U11476 ( .A(n9131), .B(n9130), .C(n15145), .D(n9129), .Z(
        n9134) );
  HS65_LL_NAND4ABX3 U11477 ( .A(n9135), .B(n9134), .C(n9133), .D(n9132), .Z(
        n9136) );
  HS65_LL_MX41X4 U11478 ( .D0(n9139), .S0(n15186), .D1(n9138), .S1(n15184), 
        .D2(n9137), .S2(n15182), .D3(n9136), .S3(n15180), .Z(n15568) );
  HS65_LLS_XOR3X2 U11479 ( .A(w2[4]), .B(n15624), .C(n15568), .Z(n9140) );
  HS65_LLS_XOR3X2 U11480 ( .A(n15583), .B(n14847), .C(n9140), .Z(n9141) );
  HS65_LL_MUX31X4 U11481 ( .D0(w2[4]), .D1(n15507), .D2(n9141), .S0(
        text_in_r[36]), .S1(n14808), .Z(N102) );
  HS65_LL_AOI12X2 U11482 ( .A(\u0/r0/rcnt [0]), .B(\u0/r0/rcnt [1]), .C(
        \u0/r0/rcnt [2]), .Z(n14988) );
  HS65_LL_NOR2X2 U11483 ( .A(n14988), .B(\u0/r0/N70 ), .Z(\u0/r0/N80 ) );
  HS65_LL_NAND2X2 U11484 ( .A(\u0/r0/rcnt [0]), .B(\u0/r0/rcnt [1]), .Z(n9142)
         );
  HS65_LL_OAI21X2 U11485 ( .A(\u0/r0/rcnt [0]), .B(\u0/r0/rcnt [1]), .C(n9142), 
        .Z(n14996) );
  HS65_LL_NOR2X2 U11486 ( .A(n15842), .B(n14996), .Z(\u0/r0/N79 ) );
  HS65_LL_IVX2 U11487 ( .A(dcnt[3]), .Z(n7664) );
  HS65_LL_IVX2 U11488 ( .A(dcnt[0]), .Z(n7668) );
  HS65_LL_IVX2 U11489 ( .A(dcnt[1]), .Z(n7665) );
  HS65_LL_NOR2X2 U11490 ( .A(n15842), .B(n14990), .Z(\u0/r0/N81 ) );
  HS65_LL_IVX2 U11491 ( .A(w3[9]), .Z(n15433) );
  HS65_LL_IVX2 U11492 ( .A(w3[14]), .Z(n15711) );
  HS65_LL_NOR2X2 U11493 ( .A(n15433), .B(n15711), .Z(n9192) );
  HS65_LL_NAND2X2 U11494 ( .A(w3[15]), .B(n9192), .Z(n9170) );
  HS65_LL_IVX2 U11495 ( .A(w3[11]), .Z(n15431) );
  HS65_LL_NAND2X2 U11496 ( .A(w3[8]), .B(n15431), .Z(n9151) );
  HS65_LL_NOR2X2 U11497 ( .A(w3[13]), .B(n9151), .Z(n9168) );
  HS65_LL_IVX2 U11498 ( .A(n9168), .Z(n9147) );
  HS65_LL_NOR2X2 U11499 ( .A(n9170), .B(n9147), .Z(n9886) );
  HS65_LL_NAND2X2 U11500 ( .A(w3[8]), .B(w3[11]), .Z(n9143) );
  HS65_LL_IVX2 U11501 ( .A(w3[15]), .Z(n15427) );
  HS65_LL_NAND2X2 U11502 ( .A(n15433), .B(n15711), .Z(n9167) );
  HS65_LL_NOR2X2 U11503 ( .A(n15427), .B(n9167), .Z(n9181) );
  HS65_LL_IVX2 U11504 ( .A(n9181), .Z(n9158) );
  HS65_LL_OR2X4 U11505 ( .A(n9143), .B(n9158), .Z(n9551) );
  HS65_LL_NOR2X2 U11506 ( .A(w3[13]), .B(n9551), .Z(n9299) );
  HS65_LL_NAND3X2 U11507 ( .A(w3[8]), .B(w3[11]), .C(w3[13]), .Z(n9198) );
  HS65_LL_NOR2X2 U11508 ( .A(n9167), .B(w3[15]), .Z(n9145) );
  HS65_LL_IVX2 U11509 ( .A(n9145), .Z(n9176) );
  HS65_LL_NOR2X2 U11510 ( .A(n9198), .B(n9176), .Z(n9550) );
  HS65_LL_IVX2 U11511 ( .A(n9550), .Z(n9317) );
  HS65_LL_NAND2AX4 U11512 ( .A(n9299), .B(n9317), .Z(n9213) );
  HS65_LL_IVX2 U11513 ( .A(n9198), .Z(n9221) );
  HS65_LL_NAND2X2 U11514 ( .A(w3[14]), .B(n15433), .Z(n9144) );
  HS65_LL_IVX2 U11515 ( .A(n9144), .Z(n9220) );
  HS65_LL_NAND2X2 U11516 ( .A(n9220), .B(n15427), .Z(n9288) );
  HS65_LL_IVX2 U11517 ( .A(n9288), .Z(n9169) );
  HS65_LL_NAND2X2 U11518 ( .A(n9221), .B(n9169), .Z(n9546) );
  HS65_LL_NOR3X1 U11519 ( .A(w3[8]), .B(w3[11]), .C(w3[13]), .Z(n9207) );
  HS65_LL_NAND2X2 U11520 ( .A(n9145), .B(n9207), .Z(n9760) );
  HS65_LL_NAND2X2 U11521 ( .A(n9546), .B(n9760), .Z(n9298) );
  HS65_LL_NAND2X2 U11522 ( .A(n15427), .B(n9192), .Z(n9228) );
  HS65_LL_IVX2 U11523 ( .A(n9228), .Z(n9157) );
  HS65_LL_NAND2X2 U11524 ( .A(n9221), .B(n9157), .Z(n9308) );
  HS65_LL_NOR2X2 U11525 ( .A(n15427), .B(n9144), .Z(n9172) );
  HS65_LL_NAND2X2 U11526 ( .A(n9172), .B(n9168), .Z(n9347) );
  HS65_LL_NAND3AX3 U11527 ( .A(n9298), .B(n9308), .C(n9347), .Z(n9757) );
  HS65_LL_NOR2X2 U11528 ( .A(n9198), .B(n9170), .Z(n9540) );
  HS65_LL_NOR2X2 U11529 ( .A(w3[8]), .B(n15431), .Z(n9156) );
  HS65_LL_NAND2X2 U11530 ( .A(n9156), .B(n15707), .Z(n9180) );
  HS65_LL_NOR2X2 U11531 ( .A(n9144), .B(n9180), .Z(n9183) );
  HS65_LL_NAND2X2 U11532 ( .A(w3[15]), .B(n9183), .Z(n9532) );
  HS65_LL_NAND2AX4 U11533 ( .A(n9540), .B(n9532), .Z(n9879) );
  HS65_LL_NAND3X2 U11534 ( .A(w3[11]), .B(w3[8]), .C(n15707), .Z(n10238) );
  HS65_LL_IVX2 U11535 ( .A(n10238), .Z(n9160) );
  HS65_LL_NAND2X2 U11536 ( .A(n9169), .B(n9160), .Z(n9314) );
  HS65_LL_IVX2 U11537 ( .A(n9314), .Z(n9300) );
  HS65_LL_NOR2X2 U11538 ( .A(w3[8]), .B(w3[11]), .Z(n9148) );
  HS65_LL_NAND2X2 U11539 ( .A(w3[13]), .B(n9148), .Z(n9287) );
  HS65_LL_NAND2X2 U11540 ( .A(w3[9]), .B(n15711), .Z(n9173) );
  HS65_LL_IVX2 U11541 ( .A(n9173), .Z(n9518) );
  HS65_LL_NAND2X2 U11542 ( .A(w3[15]), .B(n9518), .Z(n9152) );
  HS65_LL_NOR2X2 U11543 ( .A(n9287), .B(n9152), .Z(n9539) );
  HS65_LL_NOR2X2 U11544 ( .A(n9300), .B(n9539), .Z(n9337) );
  HS65_LL_NOR2X2 U11545 ( .A(n9180), .B(n9170), .Z(n9352) );
  HS65_LL_IVX2 U11546 ( .A(n9352), .Z(n9331) );
  HS65_LL_NAND2X2 U11547 ( .A(n9337), .B(n9331), .Z(n9219) );
  HS65_LL_IVX2 U11548 ( .A(n9207), .Z(n9150) );
  HS65_LL_NOR2X2 U11549 ( .A(n9170), .B(n9150), .Z(n9759) );
  HS65_LL_NOR2X2 U11550 ( .A(n15707), .B(n9151), .Z(n9517) );
  HS65_LL_IVX2 U11551 ( .A(n9517), .Z(n9191) );
  HS65_LL_NOR3X1 U11552 ( .A(w3[15]), .B(n9191), .C(n9173), .Z(n9558) );
  HS65_LL_AOI12X2 U11553 ( .A(n9145), .B(n9156), .C(n9558), .Z(n9307) );
  HS65_LL_NAND3X2 U11554 ( .A(w3[9]), .B(n9160), .C(n15427), .Z(n9304) );
  HS65_LL_NAND3AX3 U11555 ( .A(n9759), .B(n9307), .C(n9304), .Z(n9146) );
  HS65_LL_NOR3X1 U11556 ( .A(n9879), .B(n9219), .C(n9146), .Z(n10254) );
  HS65_LL_NOR2X2 U11557 ( .A(n9152), .B(n10238), .Z(n9336) );
  HS65_LL_NOR3X1 U11558 ( .A(n15433), .B(n15711), .C(n9287), .Z(n9297) );
  HS65_LL_NOR2AX3 U11559 ( .A(n9297), .B(w3[15]), .Z(n10242) );
  HS65_LL_NOR2X2 U11560 ( .A(n9287), .B(n9176), .Z(n9289) );
  HS65_LL_NOR3X1 U11561 ( .A(n9336), .B(n10242), .C(n9289), .Z(n9536) );
  HS65_LL_NAND4ABX3 U11562 ( .A(n9213), .B(n9757), .C(n10254), .D(n9536), .Z(
        n9154) );
  HS65_LL_NOR2X2 U11563 ( .A(n9151), .B(n9176), .Z(n9182) );
  HS65_LL_NOR2X2 U11564 ( .A(w3[15]), .B(n9173), .Z(n9161) );
  HS65_LL_NAND2X2 U11565 ( .A(n9221), .B(n9161), .Z(n9768) );
  HS65_LL_IVX2 U11566 ( .A(n9768), .Z(n9553) );
  HS65_LL_NOR2X2 U11567 ( .A(n9147), .B(n9152), .Z(n9346) );
  HS65_LL_NOR2X2 U11568 ( .A(n9180), .B(n9152), .Z(n10225) );
  HS65_LL_NOR2X2 U11569 ( .A(n9198), .B(n9152), .Z(n9775) );
  HS65_LL_NOR3X1 U11570 ( .A(n9346), .B(n10225), .C(n9775), .Z(n9366) );
  HS65_LL_NAND2X2 U11571 ( .A(n9517), .B(n9157), .Z(n9547) );
  HS65_LL_AND2X4 U11572 ( .A(n9148), .B(n9161), .Z(n9515) );
  HS65_LL_NAND2X2 U11573 ( .A(n15707), .B(n9515), .Z(n9223) );
  HS65_LL_IVX2 U11574 ( .A(n9223), .Z(n9763) );
  HS65_LL_IVX2 U11575 ( .A(n9172), .Z(n9197) );
  HS65_LL_NOR2X2 U11576 ( .A(n9197), .B(n9287), .Z(n9178) );
  HS65_LL_NOR4ABX2 U11577 ( .A(n9366), .B(n9547), .C(n9763), .D(n9178), .Z(
        n9891) );
  HS65_LL_NOR2X2 U11578 ( .A(n9287), .B(n9158), .Z(n9900) );
  HS65_LL_AOI12X2 U11579 ( .A(n9517), .B(n9220), .C(n9900), .Z(n9212) );
  HS65_LL_NAND2X2 U11580 ( .A(n9156), .B(n9161), .Z(n10232) );
  HS65_LL_NAND3X2 U11581 ( .A(n9891), .B(n9212), .C(n10232), .Z(n9149) );
  HS65_LL_NOR3X1 U11582 ( .A(n9182), .B(n9553), .C(n9149), .Z(n9755) );
  HS65_LL_NOR2X2 U11583 ( .A(n9197), .B(n9150), .Z(n9519) );
  HS65_LL_NOR2X2 U11584 ( .A(n9151), .B(n9158), .Z(n9534) );
  HS65_LL_NAND2X2 U11585 ( .A(w3[13]), .B(n9534), .Z(n9766) );
  HS65_LL_NAND2X2 U11586 ( .A(n9157), .B(n9207), .Z(n9528) );
  HS65_LL_NAND2X2 U11587 ( .A(n9766), .B(n9528), .Z(n9360) );
  HS65_LL_NAND2X2 U11588 ( .A(n9168), .B(n9161), .Z(n9751) );
  HS65_LL_IVX2 U11589 ( .A(n9152), .Z(n9208) );
  HS65_LL_NAND2X2 U11590 ( .A(w3[13]), .B(n9156), .Z(n9175) );
  HS65_LL_IVX2 U11591 ( .A(n9175), .Z(n9290) );
  HS65_LL_NAND2X2 U11592 ( .A(n9208), .B(n9290), .Z(n9171) );
  HS65_LL_NAND2X2 U11593 ( .A(n9751), .B(n9171), .Z(n9224) );
  HS65_LL_NOR3X1 U11594 ( .A(n9519), .B(n9360), .C(n9224), .Z(n9153) );
  HS65_LL_NAND4ABX3 U11595 ( .A(n9886), .B(n9154), .C(n9755), .D(n9153), .Z(
        n9189) );
  HS65_LL_NOR2X2 U11596 ( .A(w3[10]), .B(w3[12]), .Z(n10260) );
  HS65_LL_NAND2X2 U11597 ( .A(w3[13]), .B(n9515), .Z(n9774) );
  HS65_LL_NAND2X2 U11598 ( .A(n9157), .B(n9160), .Z(n9354) );
  HS65_LL_NAND3X2 U11599 ( .A(n9768), .B(n9774), .C(n9354), .Z(n10236) );
  HS65_LL_NOR2X2 U11600 ( .A(n9197), .B(n10238), .Z(n9320) );
  HS65_LL_NOR2AX3 U11601 ( .A(n9546), .B(n9320), .Z(n9202) );
  HS65_LL_NOR2AX3 U11602 ( .A(n9202), .B(n9519), .Z(n9340) );
  HS65_LL_IVX2 U11603 ( .A(n9340), .Z(n9913) );
  HS65_LL_OR2X4 U11604 ( .A(n9170), .B(n10238), .Z(n9901) );
  HS65_LL_NAND2X2 U11605 ( .A(n9901), .B(n9171), .Z(n9217) );
  HS65_LL_OAI21X2 U11606 ( .A(n9173), .B(n9180), .C(n9308), .Z(n9914) );
  HS65_LL_NOR3X1 U11607 ( .A(n9299), .B(n9217), .C(n9914), .Z(n9155) );
  HS65_LL_NAND2X2 U11608 ( .A(n9181), .B(n9207), .Z(n9750) );
  HS65_LL_IVX2 U11609 ( .A(n9886), .Z(n9205) );
  HS65_LL_NAND3X2 U11610 ( .A(n9155), .B(n9750), .C(n9205), .Z(n9201) );
  HS65_LL_NOR2X2 U11611 ( .A(n9183), .B(n9201), .Z(n9543) );
  HS65_LL_IVX2 U11612 ( .A(n9156), .Z(n9227) );
  HS65_LL_NOR3X1 U11613 ( .A(w3[13]), .B(n9227), .C(n9228), .Z(n9555) );
  HS65_LL_IVX2 U11614 ( .A(n9751), .Z(n9349) );
  HS65_LL_NOR2X2 U11615 ( .A(n9180), .B(n9176), .Z(n9899) );
  HS65_LL_NOR2X2 U11616 ( .A(n9170), .B(n9175), .Z(n9908) );
  HS65_LL_IVX2 U11617 ( .A(n9908), .Z(n9294) );
  HS65_LL_NAND2X2 U11618 ( .A(n9157), .B(n9168), .Z(n9520) );
  HS65_LL_NAND3X2 U11619 ( .A(n9294), .B(n9520), .C(n9347), .Z(n9177) );
  HS65_LL_NAND2X2 U11620 ( .A(n9169), .B(n9290), .Z(n9773) );
  HS65_LL_NAND2X2 U11621 ( .A(n9517), .B(n9208), .Z(n9306) );
  HS65_LL_NOR2X2 U11622 ( .A(n9158), .B(n9175), .Z(n9767) );
  HS65_LL_NOR2AX3 U11623 ( .A(n9306), .B(n9767), .Z(n10226) );
  HS65_LL_NAND4ABX3 U11624 ( .A(n9899), .B(n9177), .C(n9773), .D(n10226), .Z(
        n9159) );
  HS65_LL_NOR3X1 U11625 ( .A(n9555), .B(n9349), .C(n9159), .Z(n9895) );
  HS65_LL_NAND4ABX3 U11626 ( .A(n10236), .B(n9913), .C(n9543), .D(n9895), .Z(
        n9162) );
  HS65_LL_AND2X4 U11627 ( .A(n9161), .B(n9160), .Z(n9880) );
  HS65_LL_NOR3X1 U11628 ( .A(n9775), .B(n9880), .C(n9539), .Z(n9560) );
  HS65_LL_NAND4ABX3 U11629 ( .A(n9759), .B(n9162), .C(n9212), .D(n9560), .Z(
        n9188) );
  HS65_LL_IVX2 U11630 ( .A(w3[10]), .Z(n11559) );
  HS65_LL_NAND2X2 U11631 ( .A(w3[12]), .B(n11559), .Z(n10255) );
  HS65_LL_IVX2 U11632 ( .A(n10255), .Z(n9919) );
  HS65_LL_NOR2X2 U11633 ( .A(n15707), .B(n9551), .Z(n9319) );
  HS65_LL_NOR3X1 U11634 ( .A(w3[15]), .B(n9167), .C(n10238), .Z(n9530) );
  HS65_LL_NOR2X2 U11635 ( .A(n9759), .B(n9530), .Z(n9218) );
  HS65_LL_NAND2AX4 U11636 ( .A(n9319), .B(n9218), .Z(n9203) );
  HS65_LL_NOR2X2 U11637 ( .A(n9191), .B(n9197), .Z(n9335) );
  HS65_LL_NOR2X2 U11638 ( .A(n9335), .B(n9550), .Z(n9165) );
  HS65_LL_NOR2X2 U11639 ( .A(n9228), .B(n9175), .Z(n9353) );
  HS65_LL_NOR2X2 U11640 ( .A(n9553), .B(n9353), .Z(n9164) );
  HS65_LL_NOR3X1 U11641 ( .A(w3[15]), .B(n9173), .C(n9175), .Z(n9179) );
  HS65_LL_NAND2X2 U11642 ( .A(n15707), .B(n9534), .Z(n9226) );
  HS65_LL_IVX2 U11643 ( .A(n9226), .Z(n9195) );
  HS65_LL_NAND2X2 U11644 ( .A(n9169), .B(n9207), .Z(n10239) );
  HS65_LL_NAND2X2 U11645 ( .A(n9750), .B(n10239), .Z(n10230) );
  HS65_LL_NOR3X1 U11646 ( .A(n9195), .B(n10242), .C(n10230), .Z(n9163) );
  HS65_LL_NAND3X2 U11647 ( .A(n9163), .B(n9306), .C(n9528), .Z(n9885) );
  HS65_LL_NOR4ABX2 U11648 ( .A(n9165), .B(n9164), .C(n9179), .D(n9885), .Z(
        n9166) );
  HS65_LL_OAI112X1 U11649 ( .A(n9175), .B(n9167), .C(n9166), .D(n9760), .Z(
        n9365) );
  HS65_LL_NAND2X2 U11650 ( .A(n9169), .B(n9168), .Z(n9761) );
  HS65_LL_IVX2 U11651 ( .A(n9761), .Z(n9345) );
  HS65_LL_NOR2X2 U11652 ( .A(n9178), .B(n9345), .Z(n9211) );
  HS65_LL_NOR2X2 U11653 ( .A(n9170), .B(n9191), .Z(n9888) );
  HS65_LL_IVX2 U11654 ( .A(n9171), .Z(n9305) );
  HS65_LL_NOR4ABX2 U11655 ( .A(n9546), .B(n9211), .C(n9888), .D(n9305), .Z(
        n9904) );
  HS65_LL_AND2X4 U11656 ( .A(n9547), .B(n9751), .Z(n9309) );
  HS65_LL_NAND2X2 U11657 ( .A(n9172), .B(n9290), .Z(n9322) );
  HS65_LL_NOR3X1 U11658 ( .A(w3[15]), .B(n9180), .C(n9173), .Z(n9516) );
  HS65_LL_NOR4ABX2 U11659 ( .A(n9309), .B(n9322), .C(n9908), .D(n9516), .Z(
        n9174) );
  HS65_LL_NAND4ABX3 U11660 ( .A(n9203), .B(n9365), .C(n9904), .D(n9174), .Z(
        n9187) );
  HS65_LL_NAND2X2 U11661 ( .A(w3[10]), .B(w3[12]), .Z(n10264) );
  HS65_LL_IVX2 U11662 ( .A(n10264), .Z(n9917) );
  HS65_LL_NOR2X2 U11663 ( .A(n9176), .B(n9175), .Z(n9552) );
  HS65_LL_NOR3X1 U11664 ( .A(n9763), .B(n9552), .C(n9177), .Z(n10266) );
  HS65_LL_NOR2X2 U11665 ( .A(n9178), .B(n9336), .Z(n10233) );
  HS65_LL_NOR2X2 U11666 ( .A(n9759), .B(n9179), .Z(n9199) );
  HS65_LL_NAND2X2 U11667 ( .A(w3[13]), .B(n9182), .Z(n9525) );
  HS65_LL_IVX2 U11668 ( .A(n9180), .Z(n9193) );
  HS65_LL_NAND2X2 U11669 ( .A(n9193), .B(n9181), .Z(n9756) );
  HS65_LL_NAND2X2 U11670 ( .A(n9525), .B(n9756), .Z(n9214) );
  HS65_LL_NOR4ABX2 U11671 ( .A(n10233), .B(n9199), .C(n9298), .D(n9214), .Z(
        n9363) );
  HS65_LL_NAND2X2 U11672 ( .A(n10266), .B(n9363), .Z(n9542) );
  HS65_LL_NAND2X2 U11673 ( .A(n9774), .B(n9314), .Z(n10244) );
  HS65_LL_NOR4ABX2 U11674 ( .A(n9761), .B(n9308), .C(n9305), .D(n10244), .Z(
        n9185) );
  HS65_LL_NOR2AX3 U11675 ( .A(n9182), .B(w3[13]), .Z(n9772) );
  HS65_LL_NOR2X2 U11676 ( .A(n9772), .B(n9899), .Z(n9529) );
  HS65_LL_IVX2 U11677 ( .A(n9289), .Z(n9522) );
  HS65_LL_NOR4ABX2 U11678 ( .A(n9529), .B(n9522), .C(n9516), .D(n10242), .Z(
        n9361) );
  HS65_LL_NOR2AX3 U11679 ( .A(n9183), .B(w3[15]), .Z(n9889) );
  HS65_LL_NOR4ABX2 U11680 ( .A(n9560), .B(n9361), .C(n9889), .D(n9555), .Z(
        n9184) );
  HS65_LL_NAND4ABX3 U11681 ( .A(n9320), .B(n9542), .C(n9185), .D(n9184), .Z(
        n9186) );
  HS65_LL_IVX2 U11682 ( .A(w3[12]), .Z(n15429) );
  HS65_LL_NAND2X2 U11683 ( .A(w3[10]), .B(n15429), .Z(n10257) );
  HS65_LL_IVX2 U11684 ( .A(n10257), .Z(n9915) );
  HS65_LL_MX41X4 U11685 ( .D0(n9189), .S0(n10260), .D1(n9188), .S1(n9919), 
        .D2(n9187), .S2(n9917), .D3(n9186), .S3(n9915), .Z(n9190) );
  HS65_LLS_XNOR2X3 U11686 ( .A(w0[21]), .B(n9190), .Z(n15005) );
  HS65_LL_IVX4 U11687 ( .A(n15844), .Z(n15110) );
  HS65_LL_MUX21I1X3 U11688 ( .D0(n15005), .D1(key[117]), .S0(n15110), .Z(
        \u0/N63 ) );
  HS65_LL_NOR2X2 U11689 ( .A(n9191), .B(n9288), .Z(n9545) );
  HS65_LL_IVX2 U11690 ( .A(n9545), .Z(n9881) );
  HS65_LL_NAND2X2 U11691 ( .A(n9881), .B(n9294), .Z(n9310) );
  HS65_LL_AOI12X2 U11692 ( .A(n9193), .B(n9192), .C(n9310), .Z(n9194) );
  HS65_LL_NAND4ABX3 U11693 ( .A(n9346), .B(n9772), .C(n9522), .D(n9194), .Z(
        n9196) );
  HS65_LL_NOR2X2 U11694 ( .A(n9195), .B(n9552), .Z(n10240) );
  HS65_LL_NAND4ABX3 U11695 ( .A(n9336), .B(n9196), .C(n10240), .D(n9756), .Z(
        n9905) );
  HS65_LL_NAND2AX4 U11696 ( .A(n9320), .B(n9528), .Z(n10224) );
  HS65_LL_NAND2X2 U11697 ( .A(n9317), .B(n9773), .Z(n9348) );
  HS65_LL_NOR2X2 U11698 ( .A(n9763), .B(n9348), .Z(n10235) );
  HS65_LL_NAND4ABX3 U11699 ( .A(n9905), .B(n10224), .C(n9525), .D(n10235), .Z(
        n9200) );
  HS65_LL_NOR2X2 U11700 ( .A(n9198), .B(n9197), .Z(n9894) );
  HS65_LL_NOR2X2 U11701 ( .A(n9894), .B(n9558), .Z(n9357) );
  HS65_LL_NAND4ABX3 U11702 ( .A(n9201), .B(n9200), .C(n9199), .D(n9357), .Z(
        n9236) );
  HS65_LL_NAND4ABX3 U11703 ( .A(n9880), .B(n9203), .C(n9202), .D(n9522), .Z(
        n9204) );
  HS65_LL_NOR2X2 U11704 ( .A(n9540), .B(n9299), .Z(n9896) );
  HS65_LL_NAND4ABX3 U11705 ( .A(n9888), .B(n9204), .C(n9896), .D(n9525), .Z(
        n10237) );
  HS65_LL_NAND3AX3 U11706 ( .A(n9346), .B(n9547), .C(n9205), .Z(n9206) );
  HS65_LL_NOR3X1 U11707 ( .A(n9539), .B(n10237), .C(n9206), .Z(n9231) );
  HS65_LL_NOR3X1 U11708 ( .A(n9352), .B(n9552), .C(n9305), .Z(n9209) );
  HS65_LL_NAND2X2 U11709 ( .A(n9208), .B(n9207), .Z(n9890) );
  HS65_LL_NAND2X2 U11710 ( .A(n9890), .B(n9756), .Z(n9225) );
  HS65_LL_NOR4ABX2 U11711 ( .A(n10233), .B(n9209), .C(n9900), .D(n9225), .Z(
        n9210) );
  HS65_LL_NAND3X2 U11712 ( .A(n9895), .B(n9231), .C(n9210), .Z(n9235) );
  HS65_LL_IVX2 U11713 ( .A(n9899), .Z(n9323) );
  HS65_LL_NAND3X2 U11714 ( .A(n9223), .B(n9766), .C(n9323), .Z(n9344) );
  HS65_LL_NAND4ABX3 U11715 ( .A(n9879), .B(n9213), .C(n9212), .D(n9211), .Z(
        n9907) );
  HS65_LL_NOR3X1 U11716 ( .A(n10236), .B(n9214), .C(n9907), .Z(n9216) );
  HS65_LL_IVX2 U11717 ( .A(n9767), .Z(n9215) );
  HS65_LL_NAND3X2 U11718 ( .A(n9216), .B(n9547), .C(n9215), .Z(n9291) );
  HS65_LL_NOR2AX3 U11719 ( .A(n9218), .B(n9217), .Z(n9350) );
  HS65_LL_AOI112X2 U11720 ( .A(n9221), .B(n9220), .C(n9886), .D(n9219), .Z(
        n9222) );
  HS65_LL_NAND4ABX3 U11721 ( .A(n9344), .B(n9291), .C(n9350), .D(n9222), .Z(
        n9234) );
  HS65_LL_NAND3X2 U11722 ( .A(n9223), .B(n9750), .C(n9322), .Z(n9526) );
  HS65_LL_NOR3X1 U11723 ( .A(n9526), .B(n9225), .C(n9224), .Z(n9777) );
  HS65_LL_NAND2X2 U11724 ( .A(w3[15]), .B(n9297), .Z(n9887) );
  HS65_LL_NAND2X2 U11725 ( .A(n9226), .B(n9887), .Z(n10252) );
  HS65_LL_OAI112X1 U11726 ( .A(n9228), .B(n9227), .C(n9357), .D(n9761), .Z(
        n9229) );
  HS65_LL_NOR4ABX2 U11727 ( .A(n9323), .B(n9766), .C(n10252), .D(n9229), .Z(
        n9302) );
  HS65_LL_NAND4ABX3 U11728 ( .A(n9545), .B(n9519), .C(n9306), .D(n9347), .Z(
        n9230) );
  HS65_LL_NOR3AX2 U11729 ( .A(n9231), .B(n10236), .C(n9230), .Z(n9232) );
  HS65_LL_NAND3X2 U11730 ( .A(n9777), .B(n9302), .C(n9232), .Z(n9233) );
  HS65_LL_MX41X4 U11731 ( .D0(n9236), .S0(n10260), .D1(n9235), .S1(n9919), 
        .D2(n9234), .S2(n9917), .D3(n9233), .S3(n9915), .Z(n9237) );
  HS65_LLS_XNOR2X3 U11732 ( .A(w0[18]), .B(n9237), .Z(n10085) );
  HS65_LL_IVX4 U11733 ( .A(n15844), .Z(n11617) );
  HS65_LL_MUX21I1X3 U11734 ( .D0(n10085), .D1(key[114]), .S0(n11617), .Z(
        \u0/N60 ) );
  HS65_LL_IVX2 U11735 ( .A(w0[11]), .Z(n15352) );
  HS65_LL_NOR3X1 U11736 ( .A(n9455), .B(n9578), .C(n9238), .Z(n9267) );
  HS65_LL_IVX2 U11737 ( .A(n9239), .Z(n9816) );
  HS65_LL_NOR2X2 U11738 ( .A(n9240), .B(n9584), .Z(n9844) );
  HS65_LL_NAND2X2 U11739 ( .A(n9844), .B(n9257), .Z(n9590) );
  HS65_LL_NOR4ABX2 U11740 ( .A(n9267), .B(n9816), .C(n9241), .D(n9590), .Z(
        n9242) );
  HS65_LL_NAND3AX3 U11741 ( .A(n9581), .B(n9242), .C(n9425), .Z(n9623) );
  HS65_LL_IVX2 U11742 ( .A(n9574), .Z(n9586) );
  HS65_LL_IVX2 U11743 ( .A(n9268), .Z(n9604) );
  HS65_LL_IVX2 U11744 ( .A(n9258), .Z(n9820) );
  HS65_LL_NAND2X2 U11745 ( .A(n9820), .B(n9273), .Z(n9376) );
  HS65_LL_NOR2X2 U11746 ( .A(n9603), .B(n9618), .Z(n9390) );
  HS65_LL_NAND4ABX3 U11747 ( .A(n9604), .B(n9376), .C(n9251), .D(n9390), .Z(
        n9243) );
  HS65_LL_AOI112X2 U11748 ( .A(n9245), .B(n9244), .C(n9586), .D(n9243), .Z(
        n9246) );
  HS65_LL_NAND3X2 U11749 ( .A(n9246), .B(n9616), .C(n9849), .Z(n9808) );
  HS65_LL_NOR4ABX2 U11750 ( .A(n9410), .B(n9405), .C(n9810), .D(n9587), .Z(
        n9442) );
  HS65_LL_IVX2 U11751 ( .A(n9619), .Z(n9835) );
  HS65_LL_NOR4ABX2 U11752 ( .A(n9247), .B(n9835), .C(n9456), .D(n9605), .Z(
        n9248) );
  HS65_LL_NAND4ABX3 U11753 ( .A(n9623), .B(n9808), .C(n9442), .D(n9248), .Z(
        n9285) );
  HS65_LL_IVX2 U11754 ( .A(n9391), .Z(n9381) );
  HS65_LL_NAND2X2 U11755 ( .A(n9381), .B(n9249), .Z(n9401) );
  HS65_LL_NOR4ABX2 U11756 ( .A(n9425), .B(n9401), .C(n9863), .D(n9375), .Z(
        n9254) );
  HS65_LL_NOR2X2 U11757 ( .A(n9250), .B(n9593), .Z(n9640) );
  HS65_LL_NAND3X2 U11758 ( .A(w3[7]), .B(n9792), .C(n9793), .Z(n9399) );
  HS65_LL_NAND2X2 U11759 ( .A(n9251), .B(n9399), .Z(n9453) );
  HS65_LL_NOR4ABX2 U11760 ( .A(n9640), .B(n9435), .C(n9252), .D(n9453), .Z(
        n9253) );
  HS65_LL_NAND3X2 U11761 ( .A(n9255), .B(n9254), .C(n9253), .Z(n9601) );
  HS65_LL_NAND4ABX3 U11762 ( .A(n9619), .B(n9276), .C(n9405), .D(n9817), .Z(
        n9256) );
  HS65_LL_NOR3X1 U11763 ( .A(n9446), .B(n9601), .C(n9256), .Z(n9433) );
  HS65_LL_NAND4ABX3 U11764 ( .A(n9258), .B(n9568), .C(n9257), .D(n9433), .Z(
        n9260) );
  HS65_LL_NOR2X2 U11765 ( .A(n9603), .B(n9587), .Z(n9384) );
  HS65_LL_NAND4ABX3 U11766 ( .A(n9634), .B(n9260), .C(n9259), .D(n9384), .Z(
        n9284) );
  HS65_LL_OAI21X2 U11767 ( .A(n15746), .B(n9852), .C(n9452), .Z(n9624) );
  HS65_LL_NOR2X2 U11768 ( .A(n9262), .B(n9261), .Z(n9645) );
  HS65_LL_NAND2X2 U11769 ( .A(n9405), .B(n9401), .Z(n9278) );
  HS65_LL_NOR4ABX2 U11770 ( .A(n9399), .B(n9409), .C(n9645), .D(n9278), .Z(
        n9265) );
  HS65_LL_NAND3X2 U11771 ( .A(n9625), .B(n9839), .C(n9263), .Z(n9575) );
  HS65_LL_NOR4ABX2 U11772 ( .A(n9265), .B(n9430), .C(n9264), .D(n9575), .Z(
        n9266) );
  HS65_LL_NAND4ABX3 U11773 ( .A(n9624), .B(n9812), .C(n9844), .D(n9266), .Z(
        n9283) );
  HS65_LL_IVX2 U11774 ( .A(n9267), .Z(n9274) );
  HS65_LL_NAND2X2 U11775 ( .A(n9268), .B(n9625), .Z(n9838) );
  HS65_LL_AND2X4 U11776 ( .A(n9383), .B(n9378), .Z(n9602) );
  HS65_LL_NAND3X2 U11777 ( .A(n9270), .B(n9602), .C(n9269), .Z(n9271) );
  HS65_LL_NOR3X1 U11778 ( .A(n9272), .B(n9624), .C(n9271), .Z(n9595) );
  HS65_LL_NAND4ABX3 U11779 ( .A(n9274), .B(n9838), .C(n9273), .D(n9595), .Z(
        n9281) );
  HS65_LL_NAND2X2 U11780 ( .A(n9439), .B(n9275), .Z(n9858) );
  HS65_LL_NOR4ABX2 U11781 ( .A(n9277), .B(n9798), .C(n9276), .D(n9858), .Z(
        n9279) );
  HS65_LL_NAND2X2 U11782 ( .A(n9799), .B(n9396), .Z(n9842) );
  HS65_LL_NOR4ABX2 U11783 ( .A(n9279), .B(n9616), .C(n9842), .D(n9278), .Z(
        n9633) );
  HS65_LL_NAND4ABX3 U11784 ( .A(n9393), .B(n9281), .C(n9280), .D(n9633), .Z(
        n9282) );
  HS65_LL_MX41X4 U11785 ( .D0(n9285), .S0(n9599), .D1(n9284), .S1(n9873), .D2(
        n9283), .S2(n9609), .D3(n9282), .S3(n9461), .Z(n9286) );
  HS65_LL_MUXI21X2 U11786 ( .D0(w0[11]), .D1(n15352), .S0(n9286), .Z(n15009)
         );
  HS65_LL_MUX21I1X3 U11787 ( .D0(n15009), .D1(key[107]), .S0(n15783), .Z(
        \u0/N53 ) );
  HS65_LL_NOR2X2 U11788 ( .A(n9288), .B(n9287), .Z(n9531) );
  HS65_LL_NOR3X1 U11789 ( .A(n9531), .B(n9555), .C(n9319), .Z(n9332) );
  HS65_LL_NAND2X2 U11790 ( .A(n9332), .B(n9340), .Z(n9356) );
  HS65_LL_NOR2X2 U11791 ( .A(n9346), .B(n9289), .Z(n9296) );
  HS65_LL_NAND2X2 U11792 ( .A(n9518), .B(n9290), .Z(n9293) );
  HS65_LL_NAND2X2 U11793 ( .A(n9750), .B(n9322), .Z(n9292) );
  HS65_LL_NOR4ABX2 U11794 ( .A(n9294), .B(n9293), .C(n9292), .D(n9291), .Z(
        n9295) );
  HS65_LL_NAND4ABX3 U11795 ( .A(n9297), .B(n9356), .C(n9296), .D(n9295), .Z(
        n9328) );
  HS65_LL_NAND2X2 U11796 ( .A(n9773), .B(n9520), .Z(n9358) );
  HS65_LL_NOR3X1 U11797 ( .A(n9299), .B(n9298), .C(n9358), .Z(n9301) );
  HS65_LL_NOR4ABX2 U11798 ( .A(n9302), .B(n9301), .C(n9300), .D(n9880), .Z(
        n9303) );
  HS65_LL_NAND3X2 U11799 ( .A(n9755), .B(n9350), .C(n9303), .Z(n9327) );
  HS65_LL_IVX2 U11800 ( .A(n9353), .Z(n9538) );
  HS65_LL_NAND3X2 U11801 ( .A(n9538), .B(n9304), .C(n9766), .Z(n9898) );
  HS65_LL_NOR2X2 U11802 ( .A(n9346), .B(n9305), .Z(n9884) );
  HS65_LL_IVX2 U11803 ( .A(n9531), .Z(n9537) );
  HS65_LL_NAND2X2 U11804 ( .A(n9537), .B(n9306), .Z(n10250) );
  HS65_LL_NOR4ABX2 U11805 ( .A(n9307), .B(n9528), .C(n9530), .D(n10250), .Z(
        n9780) );
  HS65_LL_NAND3X2 U11806 ( .A(n9884), .B(n9780), .C(n9532), .Z(n9313) );
  HS65_LL_NOR3X1 U11807 ( .A(n9335), .B(n9900), .C(n9320), .Z(n10253) );
  HS65_LL_NAND2X2 U11808 ( .A(n9309), .B(n9308), .Z(n9333) );
  HS65_LL_NAND2X2 U11809 ( .A(n9901), .B(n9322), .Z(n9342) );
  HS65_LL_NOR3X1 U11810 ( .A(n9333), .B(n9310), .C(n9342), .Z(n9311) );
  HS65_LL_NAND3X2 U11811 ( .A(n9311), .B(n9761), .C(n9890), .Z(n10262) );
  HS65_LL_NOR2AX3 U11812 ( .A(n9363), .B(n10262), .Z(n9312) );
  HS65_LL_NAND4ABX3 U11813 ( .A(n9898), .B(n9313), .C(n10253), .D(n9312), .Z(
        n9326) );
  HS65_LL_NOR2X2 U11814 ( .A(n9352), .B(n9353), .Z(n9910) );
  HS65_LL_NAND2X2 U11815 ( .A(n9314), .B(n9760), .Z(n10231) );
  HS65_LL_NOR2X2 U11816 ( .A(n9886), .B(n10231), .Z(n9778) );
  HS65_LL_IVX2 U11817 ( .A(n9516), .Z(n9315) );
  HS65_LL_NAND3X2 U11818 ( .A(n9778), .B(n9774), .C(n9315), .Z(n9316) );
  HS65_LL_NOR4ABX2 U11819 ( .A(n9910), .B(n9347), .C(n9540), .D(n9316), .Z(
        n9556) );
  HS65_LL_NAND4ABX3 U11820 ( .A(n9335), .B(n9558), .C(n9354), .D(n9317), .Z(
        n9318) );
  HS65_LL_NOR3X1 U11821 ( .A(n9319), .B(n10252), .C(n9318), .Z(n9544) );
  HS65_LL_NOR2X2 U11822 ( .A(n9320), .B(n9767), .Z(n9752) );
  HS65_LL_IVX2 U11823 ( .A(n9520), .Z(n9334) );
  HS65_LL_NOR2X2 U11824 ( .A(n9888), .B(n9334), .Z(n10247) );
  HS65_LL_NAND3X2 U11825 ( .A(n9752), .B(n10247), .C(n9350), .Z(n9321) );
  HS65_LL_NOR4ABX2 U11826 ( .A(n9323), .B(n9322), .C(n9333), .D(n9321), .Z(
        n9324) );
  HS65_LL_NAND3X2 U11827 ( .A(n9556), .B(n9544), .C(n9324), .Z(n9325) );
  HS65_LL_MX41X4 U11828 ( .D0(n9328), .S0(n10260), .D1(n9327), .S1(n9919), 
        .D2(n9326), .S2(n9917), .D3(n9325), .S3(n9915), .Z(n9329) );
  HS65_LLS_XNOR2X3 U11829 ( .A(w0[23]), .B(n9329), .Z(n15007) );
  HS65_LL_MUX21I1X3 U11830 ( .D0(n15007), .D1(key[119]), .S0(n15110), .Z(
        \u0/N65 ) );
  HS65_LL_IVX2 U11831 ( .A(w0[20]), .Z(n15255) );
  HS65_LL_IVX2 U11832 ( .A(n9890), .Z(n9557) );
  HS65_LL_NOR2X2 U11833 ( .A(n9557), .B(n9888), .Z(n9330) );
  HS65_LL_NAND4ABX3 U11834 ( .A(n9552), .B(n10236), .C(n9330), .D(n9522), .Z(
        n9343) );
  HS65_LL_NAND2X2 U11835 ( .A(n9332), .B(n9331), .Z(n9364) );
  HS65_LL_NOR2X2 U11836 ( .A(n9889), .B(n9364), .Z(n9754) );
  HS65_LL_NOR3X1 U11837 ( .A(n9335), .B(n9334), .C(n9333), .Z(n9339) );
  HS65_LL_OR2X4 U11838 ( .A(n9336), .B(n9894), .Z(n9771) );
  HS65_LL_NOR4ABX2 U11839 ( .A(n9337), .B(n9887), .C(n9772), .D(n9771), .Z(
        n9338) );
  HS65_LL_NAND3X2 U11840 ( .A(n9340), .B(n9339), .C(n9338), .Z(n9762) );
  HS65_LL_NAND3AX3 U11841 ( .A(n10225), .B(n9525), .C(n9347), .Z(n9341) );
  HS65_LL_NOR3X1 U11842 ( .A(n9342), .B(n9762), .C(n9341), .Z(n9882) );
  HS65_LL_NAND4ABX3 U11843 ( .A(n9344), .B(n9343), .C(n9754), .D(n9882), .Z(
        n9372) );
  HS65_LL_NOR2X2 U11844 ( .A(n9346), .B(n9345), .Z(n9533) );
  HS65_LL_NAND4ABX3 U11845 ( .A(n9349), .B(n9348), .C(n9533), .D(n9347), .Z(
        n9351) );
  HS65_LL_NAND4ABX3 U11846 ( .A(n9352), .B(n9351), .C(n9350), .D(n10239), .Z(
        n9355) );
  HS65_LL_NOR2X2 U11847 ( .A(n9353), .B(n9771), .Z(n10245) );
  HS65_LL_NOR2X2 U11848 ( .A(n10225), .B(n9539), .Z(n9523) );
  HS65_LL_AND2X4 U11849 ( .A(n9523), .B(n9354), .Z(n9902) );
  HS65_LL_NAND4ABX3 U11850 ( .A(n9356), .B(n9355), .C(n10245), .D(n9902), .Z(
        n9371) );
  HS65_LL_NAND4ABX3 U11851 ( .A(n9553), .B(n9358), .C(n9538), .D(n9357), .Z(
        n9359) );
  HS65_LL_NOR4ABX2 U11852 ( .A(n9896), .B(n9361), .C(n9360), .D(n9359), .Z(
        n9362) );
  HS65_LL_NAND4ABX3 U11853 ( .A(n9364), .B(n10262), .C(n9363), .D(n9362), .Z(
        n9370) );
  HS65_LL_IVX2 U11854 ( .A(n9773), .Z(n9758) );
  HS65_LL_NOR2X2 U11855 ( .A(n9758), .B(n9899), .Z(n9368) );
  HS65_LL_NOR4ABX2 U11856 ( .A(n9366), .B(n9774), .C(n9771), .D(n9365), .Z(
        n9367) );
  HS65_LL_NAND4ABX3 U11857 ( .A(n9519), .B(n10237), .C(n9368), .D(n9367), .Z(
        n9369) );
  HS65_LL_MX41X4 U11858 ( .D0(n9372), .S0(n10260), .D1(n9371), .S1(n9919), 
        .D2(n9370), .S2(n9917), .D3(n9369), .S3(n9915), .Z(n9373) );
  HS65_LL_MUXI21X2 U11859 ( .D0(w0[20]), .D1(n15255), .S0(n9373), .Z(n15011)
         );
  HS65_LL_MUX21I1X3 U11860 ( .D0(n15011), .D1(key[116]), .S0(n15110), .Z(
        \u0/N62 ) );
  HS65_LL_IVX2 U11861 ( .A(w0[15]), .Z(n11348) );
  HS65_LL_NOR2X2 U11862 ( .A(n9375), .B(n9374), .Z(n9416) );
  HS65_LL_NOR3X1 U11863 ( .A(n9377), .B(n9645), .C(n9376), .Z(n9379) );
  HS65_LL_NAND3X2 U11864 ( .A(n9416), .B(n9379), .C(n9378), .Z(n9847) );
  HS65_LL_NAND2X2 U11865 ( .A(n9381), .B(n9380), .Z(n9864) );
  HS65_LL_NAND4ABX3 U11866 ( .A(n9791), .B(n9836), .C(n9382), .D(n9864), .Z(
        n9592) );
  HS65_LL_NOR2X2 U11867 ( .A(n9605), .B(n9447), .Z(n9861) );
  HS65_LL_NAND3X2 U11868 ( .A(n9861), .B(n9384), .C(n9383), .Z(n9385) );
  HS65_LL_NOR3X1 U11869 ( .A(n9863), .B(n9592), .C(n9385), .Z(n9386) );
  HS65_LL_NAND4ABX3 U11870 ( .A(n9847), .B(n9575), .C(n9631), .D(n9386), .Z(
        n9422) );
  HS65_LL_NAND3X2 U11871 ( .A(n9411), .B(n9864), .C(n9616), .Z(n9424) );
  HS65_LL_IVX2 U11872 ( .A(n9577), .Z(n9607) );
  HS65_LL_NAND3X2 U11873 ( .A(n9595), .B(n9387), .C(n9607), .Z(n9388) );
  HS65_LL_NOR3X1 U11874 ( .A(n9819), .B(n9389), .C(n9388), .Z(n9830) );
  HS65_LL_OAI112X1 U11875 ( .A(n9392), .B(n9391), .C(n9830), .D(n9390), .Z(
        n9398) );
  HS65_LL_CBI4I6X2 U11876 ( .A(w3[7]), .B(n9395), .C(n9394), .D(n9393), .Z(
        n9397) );
  HS65_LL_NAND4ABX3 U11877 ( .A(n9424), .B(n9398), .C(n9397), .D(n9396), .Z(
        n9421) );
  HS65_LL_IVX2 U11878 ( .A(n9399), .Z(n9802) );
  HS65_LL_NAND2X2 U11879 ( .A(n9625), .B(n9839), .Z(n9400) );
  HS65_LL_NOR3X1 U11880 ( .A(n9802), .B(n9801), .C(n9400), .Z(n9429) );
  HS65_LL_OAI21X2 U11881 ( .A(w3[5]), .B(n9402), .C(n9401), .Z(n9862) );
  HS65_LL_NOR4ABX2 U11882 ( .A(n9429), .B(n9403), .C(n9456), .D(n9862), .Z(
        n9823) );
  HS65_LL_NOR2X2 U11883 ( .A(n9639), .B(n9634), .Z(n9448) );
  HS65_LL_IVX2 U11884 ( .A(n9591), .Z(n9457) );
  HS65_LL_NAND2X2 U11885 ( .A(n9425), .B(n9457), .Z(n9406) );
  HS65_LL_NAND3X2 U11886 ( .A(n9449), .B(n9405), .C(n9404), .Z(n9418) );
  HS65_LL_NOR4ABX2 U11887 ( .A(n9448), .B(n9844), .C(n9406), .D(n9418), .Z(
        n9407) );
  HS65_LL_NAND3X2 U11888 ( .A(n9823), .B(n9408), .C(n9407), .Z(n9420) );
  HS65_LL_NAND2X2 U11889 ( .A(n9425), .B(n9409), .Z(n9859) );
  HS65_LL_NAND4ABX3 U11890 ( .A(n9801), .B(n9862), .C(n9411), .D(n9410), .Z(
        n9412) );
  HS65_LL_NOR3X1 U11891 ( .A(n9863), .B(n9638), .C(n9412), .Z(n9629) );
  HS65_LL_NOR2X2 U11892 ( .A(n9447), .B(n9577), .Z(n9834) );
  HS65_LL_NOR4ABX2 U11893 ( .A(n9414), .B(n9413), .C(n9838), .D(n9590), .Z(
        n9415) );
  HS65_LL_NAND3X2 U11894 ( .A(n9415), .B(n9452), .C(n9817), .Z(n9644) );
  HS65_LL_NOR4ABX2 U11895 ( .A(n9416), .B(n9834), .C(n9456), .D(n9644), .Z(
        n9417) );
  HS65_LL_NAND4ABX3 U11896 ( .A(n9859), .B(n9418), .C(n9629), .D(n9417), .Z(
        n9419) );
  HS65_LL_MX41X4 U11897 ( .D0(n9422), .S0(n9599), .D1(n9421), .S1(n9873), .D2(
        n9420), .S2(n9609), .D3(n9419), .S3(n9461), .Z(n9423) );
  HS65_LL_MUXI21X2 U11898 ( .D0(w0[15]), .D1(n11348), .S0(n9423), .Z(n15013)
         );
  HS65_LL_MUX21I1X3 U11899 ( .D0(n15013), .D1(key[111]), .S0(n11617), .Z(
        \u0/N57 ) );
  HS65_LL_IVX2 U11900 ( .A(w0[12]), .Z(n15350) );
  HS65_LL_NOR2X2 U11901 ( .A(n9604), .B(n9424), .Z(n9443) );
  HS65_LL_NOR4ABX2 U11902 ( .A(n9798), .B(n9425), .C(n9591), .D(n9624), .Z(
        n9426) );
  HS65_LL_NOR4ABX2 U11903 ( .A(n9427), .B(n9426), .C(n9579), .D(n9847), .Z(
        n9428) );
  HS65_LL_NAND3X2 U11904 ( .A(n9443), .B(n9429), .C(n9428), .Z(n9465) );
  HS65_LL_NAND2AX4 U11905 ( .A(n9456), .B(n9839), .Z(n9794) );
  HS65_LL_NOR2X2 U11906 ( .A(n9645), .B(n9450), .Z(n9431) );
  HS65_LL_NAND2X2 U11907 ( .A(n9443), .B(n9430), .Z(n9571) );
  HS65_LL_NOR4ABX2 U11908 ( .A(n9832), .B(n9431), .C(n9618), .D(n9571), .Z(
        n9432) );
  HS65_LL_NAND4ABX3 U11909 ( .A(n9434), .B(n9794), .C(n9433), .D(n9432), .Z(
        n9464) );
  HS65_LL_CBI4I1X3 U11910 ( .A(n9438), .B(n9437), .C(n9436), .D(n9435), .Z(
        n9445) );
  HS65_LL_NOR2X2 U11911 ( .A(n9638), .B(n9591), .Z(n9804) );
  HS65_LL_NAND2X2 U11912 ( .A(n9804), .B(n9439), .Z(n9841) );
  HS65_LL_NAND2X2 U11913 ( .A(n9835), .B(n9817), .Z(n9441) );
  HS65_LL_NOR2X2 U11914 ( .A(n9440), .B(n9453), .Z(n9857) );
  HS65_LL_NAND4ABX3 U11915 ( .A(n9841), .B(n9441), .C(n9857), .D(n9449), .Z(
        n9444) );
  HS65_LL_NAND4ABX3 U11916 ( .A(n9445), .B(n9444), .C(n9443), .D(n9442), .Z(
        n9463) );
  HS65_LL_NOR2X2 U11917 ( .A(n9447), .B(n9446), .Z(n9800) );
  HS65_LL_NAND4ABX3 U11918 ( .A(n9450), .B(n9618), .C(n9449), .D(n9448), .Z(
        n9451) );
  HS65_LL_NOR4ABX2 U11919 ( .A(n9800), .B(n9452), .C(n9581), .D(n9451), .Z(
        n9846) );
  HS65_LL_NOR3X1 U11920 ( .A(n9455), .B(n9454), .C(n9453), .Z(n9597) );
  HS65_LL_NOR4ABX2 U11921 ( .A(n9606), .B(n9457), .C(n9619), .D(n9456), .Z(
        n9459) );
  HS65_LL_NOR4ABX2 U11922 ( .A(n9459), .B(n9816), .C(n9603), .D(n9458), .Z(
        n9460) );
  HS65_LL_NAND3X2 U11923 ( .A(n9846), .B(n9597), .C(n9460), .Z(n9462) );
  HS65_LL_MX41X4 U11924 ( .D0(n9465), .S0(n9599), .D1(n9464), .S1(n9873), .D2(
        n9463), .S2(n9609), .D3(n9462), .S3(n9461), .Z(n9466) );
  HS65_LL_MUXI21X2 U11925 ( .D0(w0[12]), .D1(n15350), .S0(n9466), .Z(n15018)
         );
  HS65_LL_MUX21I1X3 U11926 ( .D0(n15018), .D1(key[108]), .S0(n11617), .Z(
        \u0/N54 ) );
  HS65_LL_NAND2X2 U11927 ( .A(w3[27]), .B(w3[24]), .Z(n9663) );
  HS65_LL_NOR2X2 U11928 ( .A(n15242), .B(n9663), .Z(n9481) );
  HS65_LL_IVX2 U11929 ( .A(n9481), .Z(n9701) );
  HS65_LL_IVX2 U11930 ( .A(w3[31]), .Z(n15195) );
  HS65_LL_IVX2 U11931 ( .A(w3[30]), .Z(n15666) );
  HS65_LL_NAND2X2 U11932 ( .A(w3[25]), .B(n15666), .Z(n9989) );
  HS65_LL_IVX2 U11933 ( .A(n9989), .Z(n9472) );
  HS65_LL_NAND2X2 U11934 ( .A(n15195), .B(n9472), .Z(n9477) );
  HS65_LL_NOR2X2 U11935 ( .A(n9701), .B(n9477), .Z(n9981) );
  HS65_LL_IVX2 U11936 ( .A(w3[27]), .Z(n15246) );
  HS65_LL_NOR2X2 U11937 ( .A(n15246), .B(w3[24]), .Z(n9494) );
  HS65_LL_NAND2X2 U11938 ( .A(w3[29]), .B(n9494), .Z(n9478) );
  HS65_LL_NOR2X2 U11939 ( .A(n9478), .B(n9477), .Z(n9947) );
  HS65_LL_NAND3X2 U11940 ( .A(n15242), .B(n15246), .C(w3[24]), .Z(n9988) );
  HS65_LL_NOR2X2 U11941 ( .A(w3[25]), .B(w3[30]), .Z(n10010) );
  HS65_LL_NAND2X2 U11942 ( .A(w3[31]), .B(n10010), .Z(n9662) );
  HS65_LL_NOR2X2 U11943 ( .A(n9988), .B(n9662), .Z(n9673) );
  HS65_LL_NOR2X2 U11944 ( .A(n15250), .B(n15666), .Z(n10188) );
  HS65_LL_IVX2 U11945 ( .A(n10188), .Z(n9944) );
  HS65_LL_IVX2 U11946 ( .A(w3[24]), .Z(n15661) );
  HS65_LL_NAND2X2 U11947 ( .A(n15246), .B(n15661), .Z(n9487) );
  HS65_LL_NAND2AX4 U11948 ( .A(n9487), .B(w3[29]), .Z(n9942) );
  HS65_LL_NOR3X1 U11949 ( .A(w3[31]), .B(n9944), .C(n9942), .Z(n9682) );
  HS65_LL_NOR2X2 U11950 ( .A(n9673), .B(n9682), .Z(n10008) );
  HS65_LL_NOR3X1 U11951 ( .A(w3[29]), .B(w3[27]), .C(w3[24]), .Z(n9667) );
  HS65_LL_IVX2 U11952 ( .A(n9667), .Z(n9467) );
  HS65_LL_OR2X4 U11953 ( .A(n9662), .B(n9467), .Z(n9945) );
  HS65_LL_NAND2X2 U11954 ( .A(n15250), .B(w3[30]), .Z(n9990) );
  HS65_LL_NOR2X2 U11955 ( .A(n9990), .B(w3[31]), .Z(n9497) );
  HS65_LL_NAND2X2 U11956 ( .A(n9497), .B(n9667), .Z(n10007) );
  HS65_LL_NAND2X2 U11957 ( .A(n9945), .B(n10007), .Z(n10028) );
  HS65_LL_NOR3X1 U11958 ( .A(w3[31]), .B(n15250), .C(n9467), .Z(n9676) );
  HS65_LL_NAND2X2 U11959 ( .A(w3[30]), .B(n9676), .Z(n9982) );
  HS65_LL_NAND3X2 U11960 ( .A(w3[29]), .B(w3[24]), .C(n15246), .Z(n9505) );
  HS65_LL_NOR2X2 U11961 ( .A(n9505), .B(n9989), .Z(n9680) );
  HS65_LL_NAND2X2 U11962 ( .A(w3[31]), .B(n9680), .Z(n10038) );
  HS65_LL_NAND2X2 U11963 ( .A(n9982), .B(n10038), .Z(n10019) );
  HS65_LL_NOR3AX2 U11964 ( .A(n10008), .B(n10028), .C(n10019), .Z(n9468) );
  HS65_LL_IVX2 U11965 ( .A(n9468), .Z(n10216) );
  HS65_LL_IVX2 U11966 ( .A(n9478), .Z(n9469) );
  HS65_LL_NAND3X2 U11967 ( .A(n15250), .B(n15666), .C(n9469), .Z(n9490) );
  HS65_LL_NOR3X1 U11968 ( .A(w3[31]), .B(w3[25]), .C(w3[30]), .Z(n9495) );
  HS65_LL_NAND2X2 U11969 ( .A(n9667), .B(n9495), .Z(n10293) );
  HS65_LL_NAND4ABX3 U11970 ( .A(n9947), .B(n10216), .C(n9490), .D(n10293), .Z(
        n9470) );
  HS65_LL_IVX2 U11971 ( .A(n9495), .Z(n9943) );
  HS65_LL_NOR2X2 U11972 ( .A(n9701), .B(n9943), .Z(n10029) );
  HS65_LL_NOR2X2 U11973 ( .A(n15195), .B(n9990), .Z(n9496) );
  HS65_LL_IVX2 U11974 ( .A(n9496), .Z(n9486) );
  HS65_LL_NOR2X2 U11975 ( .A(n9486), .B(n9505), .Z(n9966) );
  HS65_LL_NOR2X2 U11976 ( .A(n10029), .B(n9966), .Z(n9655) );
  HS65_LL_NAND2X2 U11977 ( .A(n10188), .B(n15195), .Z(n9479) );
  HS65_LL_IVX2 U11978 ( .A(n9479), .Z(n9476) );
  HS65_LL_NAND2X2 U11979 ( .A(n9469), .B(n9476), .Z(n10205) );
  HS65_LL_NAND4ABX3 U11980 ( .A(n9981), .B(n9470), .C(n9655), .D(n10205), .Z(
        n9963) );
  HS65_LL_NOR2X2 U11981 ( .A(n9479), .B(n9505), .Z(n9708) );
  HS65_LL_NOR2X2 U11982 ( .A(n9477), .B(n9988), .Z(n9724) );
  HS65_LL_NOR2X2 U11983 ( .A(n9708), .B(n9724), .Z(n9685) );
  HS65_LL_NAND2X2 U11984 ( .A(w3[31]), .B(n10188), .Z(n9654) );
  HS65_LL_IVX2 U11985 ( .A(n9654), .Z(n9471) );
  HS65_LL_NAND2X2 U11986 ( .A(n9494), .B(n9471), .Z(n9735) );
  HS65_LL_IVX2 U11987 ( .A(n9735), .Z(n10204) );
  HS65_LL_NOR2X2 U11988 ( .A(n9486), .B(n9478), .Z(n9937) );
  HS65_LL_AOI12X2 U11989 ( .A(w3[29]), .B(n10204), .C(n9937), .Z(n9941) );
  HS65_LL_NAND2X2 U11990 ( .A(n15242), .B(n9494), .Z(n9661) );
  HS65_LL_NOR2X2 U11991 ( .A(n9477), .B(n9661), .Z(n9689) );
  HS65_LL_IVX2 U11992 ( .A(n9689), .Z(n10026) );
  HS65_LL_NAND3X2 U11993 ( .A(n9685), .B(n9941), .C(n10026), .Z(n9473) );
  HS65_LL_NOR2X2 U11994 ( .A(n9701), .B(n9662), .Z(n9950) );
  HS65_LL_NOR2X2 U11995 ( .A(w3[29]), .B(n9663), .Z(n10187) );
  HS65_LL_NAND3X2 U11996 ( .A(n10187), .B(n10010), .C(n15195), .Z(n9923) );
  HS65_LL_NAND2X2 U11997 ( .A(n9471), .B(n9667), .Z(n10278) );
  HS65_LL_NAND2X2 U11998 ( .A(n9923), .B(n10278), .Z(n9702) );
  HS65_LL_NOR2X2 U11999 ( .A(n9950), .B(n9702), .Z(n9719) );
  HS65_LL_NOR2X2 U12000 ( .A(n9654), .B(n9505), .Z(n10037) );
  HS65_LL_NAND3X2 U12001 ( .A(n15246), .B(w3[24]), .C(n9497), .Z(n9704) );
  HS65_LL_NOR2X2 U12002 ( .A(w3[29]), .B(n9704), .Z(n9729) );
  HS65_LL_NOR2X2 U12003 ( .A(n10037), .B(n9729), .Z(n10279) );
  HS65_LL_NOR2X2 U12004 ( .A(n9486), .B(n9942), .Z(n9483) );
  HS65_LL_IVX2 U12005 ( .A(n9483), .Z(n9706) );
  HS65_LL_NAND2X2 U12006 ( .A(w3[31]), .B(n9472), .Z(n9499) );
  HS65_LL_NOR2X2 U12007 ( .A(n9478), .B(n9499), .Z(n9925) );
  HS65_LL_IVX2 U12008 ( .A(n9497), .Z(n9657) );
  HS65_LL_NOR2X2 U12009 ( .A(n9701), .B(n9657), .Z(n9930) );
  HS65_LL_NOR4ABX2 U12010 ( .A(n10279), .B(n9706), .C(n9925), .D(n9930), .Z(
        n10190) );
  HS65_LL_NAND4ABX3 U12011 ( .A(n9963), .B(n9473), .C(n9719), .D(n10190), .Z(
        n9513) );
  HS65_LL_NAND2X2 U12012 ( .A(w3[26]), .B(w3[28]), .Z(n10304) );
  HS65_LL_IVX2 U12013 ( .A(n10304), .Z(n10221) );
  HS65_LL_NAND2X2 U12014 ( .A(n10187), .B(n9496), .Z(n10020) );
  HS65_LL_NOR2AX3 U12015 ( .A(n10020), .B(n9930), .Z(n9716) );
  HS65_LL_NAND2X2 U12016 ( .A(n9496), .B(n9667), .Z(n9961) );
  HS65_LL_NAND2X2 U12017 ( .A(n9716), .B(n9961), .Z(n10209) );
  HS65_LL_NOR2X2 U12018 ( .A(n15242), .B(n9704), .Z(n10212) );
  HS65_LL_NOR2X2 U12019 ( .A(n9662), .B(n9942), .Z(n10273) );
  HS65_LL_NOR2X2 U12020 ( .A(n10273), .B(n9966), .Z(n9926) );
  HS65_LL_NAND2AX4 U12021 ( .A(n10212), .B(n9926), .Z(n9504) );
  HS65_LL_NOR2X2 U12022 ( .A(n9944), .B(n9988), .Z(n9681) );
  HS65_LL_NAND2X2 U12023 ( .A(w3[31]), .B(n9681), .Z(n10288) );
  HS65_LL_IVX2 U12024 ( .A(n10187), .Z(n9474) );
  HS65_LL_NOR2X2 U12025 ( .A(n9474), .B(n9662), .Z(n9931) );
  HS65_LL_NOR2AX3 U12026 ( .A(n10288), .B(n9931), .Z(n9506) );
  HS65_LL_NOR3X1 U12027 ( .A(n15195), .B(n9944), .C(n9474), .Z(n9703) );
  HS65_LL_IVX2 U12028 ( .A(n9703), .Z(n10191) );
  HS65_LL_IVX2 U12029 ( .A(n9925), .Z(n9714) );
  HS65_LL_NAND2X2 U12030 ( .A(n10191), .B(n9714), .Z(n9475) );
  HS65_LL_NAND2X2 U12031 ( .A(n9481), .B(n9476), .Z(n10297) );
  HS65_LL_OAI21X2 U12032 ( .A(n9989), .B(n9661), .C(n10297), .Z(n10203) );
  HS65_LL_NOR4ABX2 U12033 ( .A(n9506), .B(n9945), .C(n9475), .D(n10203), .Z(
        n9743) );
  HS65_LL_OAI21X2 U12034 ( .A(n9990), .B(n9661), .C(n9743), .Z(n9658) );
  HS65_LL_NAND2X2 U12035 ( .A(n10187), .B(n9476), .Z(n9984) );
  HS65_LL_NOR2X2 U12036 ( .A(n9477), .B(n9487), .Z(n9489) );
  HS65_LL_NAND2X2 U12037 ( .A(w3[29]), .B(n9489), .Z(n9960) );
  HS65_LL_NAND2X2 U12038 ( .A(n9984), .B(n9960), .Z(n9710) );
  HS65_LL_NOR2X2 U12039 ( .A(n9981), .B(n9710), .Z(n10027) );
  HS65_LL_NAND4ABX3 U12040 ( .A(n9504), .B(n9658), .C(n10027), .D(n10278), .Z(
        n9482) );
  HS65_LL_NOR2X2 U12041 ( .A(n9486), .B(n9988), .Z(n10292) );
  HS65_LL_AOI12X2 U12042 ( .A(n10204), .B(w3[29]), .C(n10292), .Z(n9491) );
  HS65_LL_NOR2X2 U12043 ( .A(n9478), .B(n9657), .Z(n9986) );
  HS65_LL_NOR2AX3 U12044 ( .A(n9681), .B(w3[31]), .Z(n9935) );
  HS65_LL_NOR2X2 U12045 ( .A(n9986), .B(n9935), .Z(n9979) );
  HS65_LL_NOR2X2 U12046 ( .A(n9479), .B(n9661), .Z(n9948) );
  HS65_LL_NAND3X2 U12047 ( .A(n9494), .B(n9495), .C(n15242), .Z(n10182) );
  HS65_LL_IVX2 U12048 ( .A(n10182), .Z(n9973) );
  HS65_LL_NOR2X2 U12049 ( .A(n9948), .B(n9973), .Z(n9728) );
  HS65_LL_NOR2X2 U12050 ( .A(n15195), .B(n9490), .Z(n9688) );
  HS65_LL_IVX2 U12051 ( .A(n9688), .Z(n10015) );
  HS65_LL_NAND3X2 U12052 ( .A(n9979), .B(n9728), .C(n10015), .Z(n9480) );
  HS65_LL_NOR4ABX2 U12053 ( .A(n9491), .B(n10038), .C(n9724), .D(n9480), .Z(
        n10192) );
  HS65_LL_NAND3X2 U12054 ( .A(w3[25]), .B(n10187), .C(n15195), .Z(n9687) );
  HS65_LL_NOR2X2 U12055 ( .A(w3[30]), .B(n9687), .Z(n10213) );
  HS65_LL_NOR2X2 U12056 ( .A(n9499), .B(n9942), .Z(n9721) );
  HS65_LL_IVX2 U12057 ( .A(n9499), .Z(n9668) );
  HS65_LL_NAND2X2 U12058 ( .A(n9481), .B(n9668), .Z(n9959) );
  HS65_LL_IVX2 U12059 ( .A(n9959), .Z(n9679) );
  HS65_LL_NOR3X1 U12060 ( .A(n10213), .B(n9721), .C(n9679), .Z(n9671) );
  HS65_LL_NAND4ABX3 U12061 ( .A(n10209), .B(n9482), .C(n10192), .D(n9671), .Z(
        n9512) );
  HS65_LL_IVX2 U12062 ( .A(w3[28]), .Z(n15244) );
  HS65_LL_NOR2X2 U12063 ( .A(w3[26]), .B(n15244), .Z(n10308) );
  HS65_LL_NAND2X2 U12064 ( .A(n10297), .B(n9714), .Z(n9493) );
  HS65_LL_NOR2X2 U12065 ( .A(n9988), .B(n9943), .Z(n10290) );
  HS65_LL_IVX2 U12066 ( .A(n10290), .Z(n9675) );
  HS65_LL_NAND2X2 U12067 ( .A(n10026), .B(n9675), .Z(n9503) );
  HS65_LL_NAND2X2 U12068 ( .A(n10187), .B(n9668), .Z(n9958) );
  HS65_LL_IVX2 U12069 ( .A(n9958), .Z(n9674) );
  HS65_LL_NOR2X2 U12070 ( .A(n9483), .B(n9674), .Z(n10017) );
  HS65_LL_NOR2X2 U12071 ( .A(n9662), .B(n9661), .Z(n9725) );
  HS65_LL_NOR2X2 U12072 ( .A(n9930), .B(n9725), .Z(n10294) );
  HS65_LL_NOR2X2 U12073 ( .A(n9505), .B(n9943), .Z(n9715) );
  HS65_LL_NAND2AX4 U12074 ( .A(n9715), .B(n10278), .Z(n9733) );
  HS65_LL_IVX2 U12075 ( .A(n9947), .Z(n9501) );
  HS65_LL_NAND2X2 U12076 ( .A(n10293), .B(n9501), .Z(n9484) );
  HS65_LL_NOR4ABX2 U12077 ( .A(n10017), .B(n10294), .C(n9733), .D(n9484), .Z(
        n9929) );
  HS65_LL_NOR2X2 U12078 ( .A(n9942), .B(n9943), .Z(n9974) );
  HS65_LL_NOR2X2 U12079 ( .A(n9974), .B(n9973), .Z(n9485) );
  HS65_LL_NAND4ABX3 U12080 ( .A(n9682), .B(n9503), .C(n9929), .D(n9485), .Z(
        n9978) );
  HS65_LL_NOR2X2 U12081 ( .A(n9663), .B(n9486), .Z(n9734) );
  HS65_LL_OAI112X1 U12082 ( .A(n9497), .B(n9734), .C(n15242), .D(n9487), .Z(
        n9488) );
  HS65_LL_NAND4ABX3 U12083 ( .A(n9948), .B(n9978), .C(n9960), .D(n9488), .Z(
        n9492) );
  HS65_LL_IVX2 U12084 ( .A(n9489), .Z(n10041) );
  HS65_LL_NOR2X2 U12085 ( .A(w3[29]), .B(n10041), .Z(n10281) );
  HS65_LL_NOR2X2 U12086 ( .A(w3[31]), .B(n9490), .Z(n10009) );
  HS65_LL_NOR2X2 U12087 ( .A(n10281), .B(n10009), .Z(n9976) );
  HS65_LL_NAND2X2 U12088 ( .A(n9491), .B(n9976), .Z(n9660) );
  HS65_LL_NOR2X2 U12089 ( .A(n9935), .B(n9660), .Z(n10018) );
  HS65_LL_NAND4ABX3 U12090 ( .A(n9493), .B(n9492), .C(n10018), .D(n9671), .Z(
        n9511) );
  HS65_LL_IVX2 U12091 ( .A(w3[26]), .Z(n15248) );
  HS65_LL_NOR2X2 U12092 ( .A(w3[28]), .B(n15248), .Z(n10300) );
  HS65_LL_NAND2X2 U12093 ( .A(n15195), .B(n9680), .Z(n9727) );
  HS65_LL_IVX2 U12094 ( .A(n9727), .Z(n9740) );
  HS65_LL_AOI12X2 U12095 ( .A(n9495), .B(n9494), .C(n9740), .Z(n9924) );
  HS65_LL_NAND2AX4 U12096 ( .A(n9661), .B(n9496), .Z(n9927) );
  HS65_LL_NOR2X2 U12097 ( .A(n9654), .B(n9701), .Z(n9705) );
  HS65_LL_NOR2AX3 U12098 ( .A(n9927), .B(n9705), .Z(n10211) );
  HS65_LL_NAND2X2 U12099 ( .A(n10204), .B(n15242), .Z(n9970) );
  HS65_LL_IVX2 U12100 ( .A(n9970), .Z(n10272) );
  HS65_LL_NAND2X2 U12101 ( .A(n10187), .B(n9497), .Z(n10011) );
  HS65_LL_IVX2 U12102 ( .A(n9721), .Z(n10183) );
  HS65_LL_NAND2X2 U12103 ( .A(n10011), .B(n10183), .Z(n9968) );
  HS65_LL_NOR4ABX2 U12104 ( .A(n10278), .B(n9687), .C(n10272), .D(n9968), .Z(
        n9498) );
  HS65_LL_NAND3X2 U12105 ( .A(n9924), .B(n10211), .C(n9498), .Z(n10046) );
  HS65_LL_NOR3X1 U12106 ( .A(w3[25]), .B(w3[31]), .C(n9701), .Z(n9665) );
  HS65_LL_NOR2AX3 U12107 ( .A(n9961), .B(n10292), .Z(n9730) );
  HS65_LL_NAND4ABX3 U12108 ( .A(n9925), .B(n9665), .C(n9730), .D(n10297), .Z(
        n9509) );
  HS65_LL_NOR2X2 U12109 ( .A(n9499), .B(n9661), .Z(n10184) );
  HS65_LL_NOR2X2 U12110 ( .A(n9988), .B(n9499), .Z(n10270) );
  HS65_LL_NOR2X2 U12111 ( .A(n9708), .B(n10270), .Z(n9720) );
  HS65_LL_NAND3X2 U12112 ( .A(n9720), .B(n9706), .C(n9959), .Z(n9500) );
  HS65_LL_NOR3X1 U12113 ( .A(n10281), .B(n10184), .C(n9500), .Z(n10198) );
  HS65_LL_NOR2X2 U12114 ( .A(n9715), .B(n9981), .Z(n10269) );
  HS65_LL_NAND3X2 U12115 ( .A(n10198), .B(n10269), .C(n9501), .Z(n9502) );
  HS65_LL_NOR3X1 U12116 ( .A(n9504), .B(n9503), .C(n9502), .Z(n10006) );
  HS65_LL_NOR2X2 U12117 ( .A(n9505), .B(n9662), .Z(n9972) );
  HS65_LL_NOR2X2 U12118 ( .A(n9972), .B(n9682), .Z(n9678) );
  HS65_LL_NAND4ABX3 U12119 ( .A(n9974), .B(n9674), .C(n9506), .D(n9678), .Z(
        n9507) );
  HS65_LL_NOR4ABX2 U12120 ( .A(n10006), .B(n10293), .C(n9724), .D(n9507), .Z(
        n9508) );
  HS65_LL_NAND4ABX3 U12121 ( .A(n10046), .B(n9509), .C(n9508), .D(n9982), .Z(
        n9510) );
  HS65_LL_NOR2X2 U12122 ( .A(w3[26]), .B(w3[28]), .Z(n10217) );
  HS65_LL_MX41X4 U12123 ( .D0(n9513), .S0(n10221), .D1(n9512), .S1(n10308), 
        .D2(n9511), .S2(n10300), .D3(n9510), .S3(n10217), .Z(n9514) );
  HS65_LLS_XNOR2X3 U12124 ( .A(w0[5]), .B(n9514), .Z(n15016) );
  HS65_LL_MUX21I1X3 U12125 ( .D0(n15016), .D1(key[101]), .S0(n15783), .Z(
        \u0/N47 ) );
  HS65_LL_IVX2 U12126 ( .A(w0[17]), .Z(n15260) );
  HS65_LL_NOR3X1 U12127 ( .A(n9515), .B(n9894), .C(n10262), .Z(n10248) );
  HS65_LL_NOR3X1 U12128 ( .A(n9767), .B(n9516), .C(n9898), .Z(n9786) );
  HS65_LL_AOI112X2 U12129 ( .A(n9518), .B(n9517), .C(n9775), .D(n9889), .Z(
        n9909) );
  HS65_LL_NOR4ABX2 U12130 ( .A(n9551), .B(n9520), .C(n10242), .D(n9519), .Z(
        n9521) );
  HS65_LL_NAND3X2 U12131 ( .A(n9778), .B(n9909), .C(n9521), .Z(n9906) );
  HS65_LL_NOR4ABX2 U12132 ( .A(n9523), .B(n9522), .C(n9555), .D(n9906), .Z(
        n9524) );
  HS65_LL_NAND3X2 U12133 ( .A(n10248), .B(n9786), .C(n9524), .Z(n9565) );
  HS65_LL_NAND2X2 U12134 ( .A(n10239), .B(n9525), .Z(n10249) );
  HS65_LL_NAND4ABX3 U12135 ( .A(n10249), .B(n9526), .C(n9901), .D(n9887), .Z(
        n9527) );
  HS65_LL_NOR4ABX2 U12136 ( .A(n9529), .B(n9528), .C(n9555), .D(n9527), .Z(
        n9912) );
  HS65_LL_NOR4ABX2 U12137 ( .A(n9533), .B(n9532), .C(n9531), .D(n9530), .Z(
        n9770) );
  HS65_LL_NOR4ABX2 U12138 ( .A(n9912), .B(n9770), .C(n9534), .D(n9880), .Z(
        n9535) );
  HS65_LL_AOI13X2 U12139 ( .A(n9536), .B(n9556), .C(n9535), .D(n10257), .Z(
        n9564) );
  HS65_LL_NAND4ABX3 U12140 ( .A(n9540), .B(n9539), .C(n9538), .D(n9537), .Z(
        n9541) );
  HS65_LL_NOR4ABX2 U12141 ( .A(n9544), .B(n9543), .C(n9542), .D(n9541), .Z(
        n9562) );
  HS65_LL_NOR2X2 U12142 ( .A(n9545), .B(n9900), .Z(n9548) );
  HS65_LL_NAND3X2 U12143 ( .A(n9548), .B(n9547), .C(n9546), .Z(n9549) );
  HS65_LL_NOR3X1 U12144 ( .A(n9550), .B(n9772), .C(n9549), .Z(n10229) );
  HS65_LL_NAND4ABX3 U12145 ( .A(n9553), .B(n9552), .C(n9551), .D(n9756), .Z(
        n9554) );
  HS65_LL_NOR3X1 U12146 ( .A(n9889), .B(n9555), .C(n9554), .Z(n9765) );
  HS65_LL_NAND4ABX3 U12147 ( .A(n9558), .B(n9557), .C(n9556), .D(n9765), .Z(
        n9559) );
  HS65_LL_NOR4ABX2 U12148 ( .A(n10229), .B(n9560), .C(n10249), .D(n9559), .Z(
        n9561) );
  HS65_LL_OAI22X1 U12149 ( .A(n9562), .B(n10264), .C(n9561), .D(n10255), .Z(
        n9563) );
  HS65_LL_AOI112X2 U12150 ( .A(n10260), .B(n9565), .C(n9564), .D(n9563), .Z(
        n9566) );
  HS65_LL_MUXI21X2 U12151 ( .D0(n15260), .D1(w0[17]), .S0(n9566), .Z(n15020)
         );
  HS65_LL_MUX21I1X3 U12152 ( .D0(n15020), .D1(key[113]), .S0(n11617), .Z(
        \u0/N59 ) );
  HS65_LL_IVX2 U12153 ( .A(w0[14]), .Z(n15348) );
  HS65_LL_NAND4ABX3 U12154 ( .A(n9569), .B(n9568), .C(n9567), .D(n9834), .Z(
        n9570) );
  HS65_LL_NOR3X1 U12155 ( .A(n9572), .B(n9571), .C(n9570), .Z(n9856) );
  HS65_LL_NOR4ABX2 U12156 ( .A(n9856), .B(n9574), .C(n9591), .D(n9573), .Z(
        n9614) );
  HS65_LL_IVX2 U12157 ( .A(n9873), .Z(n9613) );
  HS65_LL_NOR3X1 U12158 ( .A(n9577), .B(n9576), .C(n9575), .Z(n9621) );
  HS65_LL_NAND4ABX3 U12159 ( .A(n9579), .B(n9578), .C(n9849), .D(n9616), .Z(
        n9580) );
  HS65_LL_NOR3X1 U12160 ( .A(n9581), .B(n9586), .C(n9580), .Z(n9642) );
  HS65_LL_NAND2X2 U12161 ( .A(n9799), .B(n9582), .Z(n9790) );
  HS65_LL_NOR3X1 U12162 ( .A(n9584), .B(n9790), .C(n9583), .Z(n9585) );
  HS65_LL_NAND3X2 U12163 ( .A(n9621), .B(n9642), .C(n9585), .Z(n9600) );
  HS65_LL_NOR3X1 U12164 ( .A(n9645), .B(n9587), .C(n9586), .Z(n9815) );
  HS65_LL_IVX2 U12165 ( .A(n9815), .Z(n9588) );
  HS65_LL_NOR3AX2 U12166 ( .A(n9589), .B(n9588), .C(n9842), .Z(n9821) );
  HS65_LL_NOR3X1 U12167 ( .A(n9634), .B(n9591), .C(n9590), .Z(n9594) );
  HS65_LL_NOR4ABX2 U12168 ( .A(n9595), .B(n9594), .C(n9593), .D(n9592), .Z(
        n9596) );
  HS65_LL_AOI13X2 U12169 ( .A(n9597), .B(n9821), .C(n9596), .D(n9854), .Z(
        n9598) );
  HS65_LL_CBI4I6X2 U12170 ( .A(n9601), .B(n9600), .C(n9599), .D(n9598), .Z(
        n9612) );
  HS65_LL_NAND4ABX3 U12171 ( .A(n9603), .B(n9791), .C(n9602), .D(n9864), .Z(
        n9637) );
  HS65_LL_NOR2X2 U12172 ( .A(n9605), .B(n9604), .Z(n9813) );
  HS65_LL_NAND3X2 U12173 ( .A(n9821), .B(n9813), .C(n9606), .Z(n9608) );
  HS65_LL_NAND4ABX3 U12174 ( .A(n9858), .B(n9608), .C(n9607), .D(n9839), .Z(
        n9610) );
  HS65_LL_OAI13X1 U12175 ( .A(n9623), .B(n9637), .C(n9610), .D(n9609), .Z(
        n9611) );
  HS65_LL_OAI112X1 U12176 ( .A(n9614), .B(n9613), .C(n9612), .D(n9611), .Z(
        n9615) );
  HS65_LL_MUXI21X2 U12177 ( .D0(w0[14]), .D1(n15348), .S0(n9615), .Z(n15022)
         );
  HS65_LL_MUX21I1X3 U12178 ( .D0(n15022), .D1(key[110]), .S0(n11617), .Z(
        \u0/N56 ) );
  HS65_LL_IVX2 U12179 ( .A(w0[9]), .Z(n15356) );
  HS65_LL_IVX2 U12180 ( .A(n9810), .Z(n9617) );
  HS65_LL_NAND4ABX3 U12181 ( .A(n9619), .B(n9618), .C(n9617), .D(n9616), .Z(
        n9622) );
  HS65_LL_NOR3X1 U12182 ( .A(n9802), .B(n9620), .C(n9847), .Z(n9869) );
  HS65_LL_NAND4ABX3 U12183 ( .A(n9623), .B(n9622), .C(n9869), .D(n9621), .Z(
        n9652) );
  HS65_LL_NOR4ABX2 U12184 ( .A(n9864), .B(n9625), .C(n9810), .D(n9624), .Z(
        n9628) );
  HS65_LL_NOR4ABX2 U12185 ( .A(n9629), .B(n9628), .C(n9627), .D(n9626), .Z(
        n9630) );
  HS65_LL_AOI13X2 U12186 ( .A(n9631), .B(n9840), .C(n9630), .D(n9875), .Z(
        n9651) );
  HS65_LL_NAND4ABX3 U12187 ( .A(n9635), .B(n9634), .C(n9633), .D(n9632), .Z(
        n9636) );
  HS65_LL_NOR3X1 U12188 ( .A(n9644), .B(n9637), .C(n9636), .Z(n9649) );
  HS65_LL_NOR4ABX2 U12189 ( .A(n9641), .B(n9640), .C(n9639), .D(n9638), .Z(
        n9877) );
  HS65_LL_NAND4ABX3 U12190 ( .A(n9645), .B(n9644), .C(n9643), .D(n9642), .Z(
        n9646) );
  HS65_LL_NOR4ABX2 U12191 ( .A(n9877), .B(n9647), .C(n9858), .D(n9646), .Z(
        n9648) );
  HS65_LL_OAI22X1 U12192 ( .A(n9649), .B(n9854), .C(n9648), .D(n9866), .Z(
        n9650) );
  HS65_LL_AOI112X2 U12193 ( .A(n9873), .B(n9652), .C(n9651), .D(n9650), .Z(
        n9653) );
  HS65_LL_MUXI21X2 U12194 ( .D0(n15356), .D1(w0[9]), .S0(n9653), .Z(n15030) );
  HS65_LL_MUX21I1X3 U12195 ( .D0(n15030), .D1(key[105]), .S0(n11617), .Z(
        \u0/N51 ) );
  HS65_LL_IVX2 U12196 ( .A(w0[1]), .Z(n15558) );
  HS65_LL_NOR2X2 U12197 ( .A(n9654), .B(n9942), .Z(n10202) );
  HS65_LL_NOR2X2 U12198 ( .A(n9673), .B(n10202), .Z(n10040) );
  HS65_LL_NOR4ABX2 U12199 ( .A(n9655), .B(n9984), .C(n9950), .D(n9740), .Z(
        n9656) );
  HS65_LL_NAND2X2 U12200 ( .A(n10040), .B(n9656), .Z(n9936) );
  HS65_LL_NOR2X2 U12201 ( .A(n9657), .B(n9942), .Z(n9949) );
  HS65_LL_NOR2X2 U12202 ( .A(n9935), .B(n9949), .Z(n10042) );
  HS65_LL_AND2X4 U12203 ( .A(n10205), .B(n10183), .Z(n9987) );
  HS65_LL_NOR4ABX2 U12204 ( .A(n10042), .B(n9987), .C(n9705), .D(n9658), .Z(
        n9659) );
  HS65_LL_NAND4ABX3 U12205 ( .A(n9660), .B(n9936), .C(n9929), .D(n9659), .Z(
        n9699) );
  HS65_LL_NOR2X2 U12206 ( .A(n10009), .B(n9725), .Z(n9738) );
  HS65_LL_NOR2X2 U12207 ( .A(n9981), .B(n9948), .Z(n9664) );
  HS65_LL_NOR3X1 U12208 ( .A(w3[31]), .B(n9990), .C(n9661), .Z(n10196) );
  HS65_LL_NOR2X2 U12209 ( .A(n9663), .B(n9662), .Z(n9684) );
  HS65_LL_NOR4ABX2 U12210 ( .A(n9738), .B(n9664), .C(n10196), .D(n9684), .Z(
        n10283) );
  HS65_LL_NOR2X2 U12211 ( .A(n10212), .B(n10290), .Z(n9739) );
  HS65_LL_IVX2 U12212 ( .A(n10273), .Z(n9666) );
  HS65_LL_NOR4ABX2 U12213 ( .A(n9739), .B(n9666), .C(n9708), .D(n9665), .Z(
        n10023) );
  HS65_LL_NAND2X2 U12214 ( .A(n9668), .B(n9667), .Z(n10199) );
  HS65_LL_IVX2 U12215 ( .A(n10007), .Z(n10271) );
  HS65_LL_NOR2X2 U12216 ( .A(n9715), .B(n10271), .Z(n10039) );
  HS65_LL_NAND2X2 U12217 ( .A(n10011), .B(n9970), .Z(n9669) );
  HS65_LL_NOR4ABX2 U12218 ( .A(n10293), .B(n10288), .C(n10292), .D(n9669), .Z(
        n9670) );
  HS65_LL_NAND2X2 U12219 ( .A(n9960), .B(n10205), .Z(n10014) );
  HS65_LL_NOR4ABX2 U12220 ( .A(n9670), .B(n10026), .C(n9705), .D(n10014), .Z(
        n9940) );
  HS65_LL_NAND3X2 U12221 ( .A(n10039), .B(n9671), .C(n9940), .Z(n9672) );
  HS65_LL_NOR4ABX2 U12222 ( .A(n10023), .B(n10199), .C(n9740), .D(n9672), .Z(
        n9697) );
  HS65_LL_IVX2 U12223 ( .A(n10308), .Z(n9696) );
  HS65_LL_NOR3X1 U12224 ( .A(n9674), .B(n9673), .C(n10270), .Z(n9736) );
  HS65_LL_NOR4ABX2 U12225 ( .A(n9923), .B(n9927), .C(n9949), .D(n9729), .Z(
        n10268) );
  HS65_LL_NAND3X2 U12226 ( .A(n9736), .B(n10268), .C(n9940), .Z(n9694) );
  HS65_LL_NOR2X2 U12227 ( .A(n10213), .B(n9974), .Z(n9718) );
  HS65_LL_NOR3X1 U12228 ( .A(n9703), .B(n9937), .C(n9715), .Z(n9969) );
  HS65_LL_NAND4ABX3 U12229 ( .A(n9676), .B(n10202), .C(n9728), .D(n9675), .Z(
        n9677) );
  HS65_LL_NOR3AX2 U12230 ( .A(n9969), .B(n10028), .C(n9677), .Z(n10206) );
  HS65_LL_NAND3X2 U12231 ( .A(n9718), .B(n10206), .C(n9678), .Z(n9693) );
  HS65_LL_NAND2X2 U12232 ( .A(n10293), .B(n10011), .Z(n10194) );
  HS65_LL_NOR3X1 U12233 ( .A(n9680), .B(n9679), .C(n10196), .Z(n10208) );
  HS65_LL_NAND4ABX3 U12234 ( .A(n9682), .B(n9681), .C(n9961), .D(n10208), .Z(
        n9683) );
  HS65_LL_NOR3X1 U12235 ( .A(n9684), .B(n10194), .C(n9683), .Z(n10274) );
  HS65_LL_NAND2X2 U12236 ( .A(n9685), .B(n10297), .Z(n9934) );
  HS65_LL_NAND3X2 U12237 ( .A(n9941), .B(n9704), .C(n10199), .Z(n9686) );
  HS65_LL_NOR3X1 U12238 ( .A(n9703), .B(n9934), .C(n9686), .Z(n10031) );
  HS65_LL_NOR2AX3 U12239 ( .A(n10205), .B(n9972), .Z(n10016) );
  HS65_LL_NAND2X2 U12240 ( .A(n10016), .B(n9687), .Z(n10201) );
  HS65_LL_NOR3X1 U12241 ( .A(n9689), .B(n9688), .C(n10201), .Z(n10282) );
  HS65_LL_NAND2X2 U12242 ( .A(w3[29]), .B(n9734), .Z(n10036) );
  HS65_LL_NAND4ABX3 U12243 ( .A(n10184), .B(n9948), .C(n10041), .D(n10183), 
        .Z(n9690) );
  HS65_LL_NOR4ABX2 U12244 ( .A(n10282), .B(n10036), .C(n9974), .D(n9690), .Z(
        n9691) );
  HS65_LL_IVX2 U12245 ( .A(n10217), .Z(n10295) );
  HS65_LL_AOI13X2 U12246 ( .A(n10274), .B(n10031), .C(n9691), .D(n10295), .Z(
        n9692) );
  HS65_LL_CBI4I6X2 U12247 ( .A(n9694), .B(n9693), .C(n10300), .D(n9692), .Z(
        n9695) );
  HS65_LL_CBI4I1X3 U12248 ( .A(n10283), .B(n9697), .C(n9696), .D(n9695), .Z(
        n9698) );
  HS65_LL_AOI12X2 U12249 ( .A(n10221), .B(n9699), .C(n9698), .Z(n9700) );
  HS65_LL_MUXI21X2 U12250 ( .D0(n15558), .D1(w0[1]), .S0(n9700), .Z(n15032) );
  HS65_LL_MUX21I1X3 U12251 ( .D0(n15032), .D1(key[97]), .S0(n15783), .Z(
        \u0/N43 ) );
  HS65_LL_OAI112X1 U12252 ( .A(n9701), .B(n9990), .C(n10011), .D(n9970), .Z(
        n9713) );
  HS65_LL_NOR3X1 U12253 ( .A(n9703), .B(n9925), .C(n9702), .Z(n9985) );
  HS65_LL_NAND3X2 U12254 ( .A(n9926), .B(n9704), .C(n9927), .Z(n9707) );
  HS65_LL_NOR2X2 U12255 ( .A(n9931), .B(n9705), .Z(n10197) );
  HS65_LL_NAND4ABX3 U12256 ( .A(n10029), .B(n9707), .C(n10197), .D(n9706), .Z(
        n10302) );
  HS65_LL_NAND4ABX3 U12257 ( .A(n9708), .B(n9725), .C(n10015), .D(n10269), .Z(
        n9709) );
  HS65_LL_NOR3X1 U12258 ( .A(n9710), .B(n10302), .C(n9709), .Z(n9951) );
  HS65_LL_NAND2X2 U12259 ( .A(n10183), .B(n10288), .Z(n9711) );
  HS65_LL_NOR4ABX2 U12260 ( .A(n9951), .B(n10182), .C(n10281), .D(n9711), .Z(
        n9712) );
  HS65_LL_NAND4ABX3 U12261 ( .A(n9972), .B(n9713), .C(n9985), .D(n9712), .Z(
        n9747) );
  HS65_LL_IVX2 U12262 ( .A(n10017), .Z(n10032) );
  HS65_LL_NAND2X2 U12263 ( .A(n10199), .B(n9714), .Z(n9723) );
  HS65_LL_NOR4ABX2 U12264 ( .A(n10197), .B(n9716), .C(n9715), .D(n10037), .Z(
        n9717) );
  HS65_LL_NAND3X2 U12265 ( .A(n9719), .B(n9718), .C(n9717), .Z(n10034) );
  HS65_LL_NAND4ABX3 U12266 ( .A(n9721), .B(n10034), .C(n9720), .D(n10288), .Z(
        n9732) );
  HS65_LL_NOR4ABX2 U12267 ( .A(n9970), .B(n9738), .C(n10273), .D(n9732), .Z(
        n9722) );
  HS65_LL_NAND4ABX3 U12268 ( .A(n10032), .B(n9723), .C(n10192), .D(n9722), .Z(
        n9746) );
  HS65_LL_NAND2AX4 U12269 ( .A(n9724), .B(n9945), .Z(n10002) );
  HS65_LL_NOR3X1 U12270 ( .A(n9937), .B(n9725), .C(n10002), .Z(n9726) );
  HS65_LL_NAND4ABX3 U12271 ( .A(n10281), .B(n9925), .C(n9726), .D(n10199), .Z(
        n10310) );
  HS65_LL_NAND3X2 U12272 ( .A(n10016), .B(n9727), .C(n10036), .Z(n9980) );
  HS65_LL_NAND4ABX3 U12273 ( .A(n9729), .B(n9980), .C(n9728), .D(n10040), .Z(
        n9933) );
  HS65_LL_NOR4ABX2 U12274 ( .A(n9730), .B(n10038), .C(n10212), .D(n9933), .Z(
        n9731) );
  HS65_LL_NAND4ABX3 U12275 ( .A(n9732), .B(n10310), .C(n10027), .D(n9731), .Z(
        n9745) );
  HS65_LL_NOR3X1 U12276 ( .A(n10029), .B(n9734), .C(n9733), .Z(n9742) );
  HS65_LL_NOR3X1 U12277 ( .A(n9947), .B(n10281), .C(n9986), .Z(n10030) );
  HS65_LL_NOR4ABX2 U12278 ( .A(n9736), .B(n9735), .C(n9974), .D(n9948), .Z(
        n9737) );
  HS65_LL_NAND3X2 U12279 ( .A(n9739), .B(n9738), .C(n9737), .Z(n10186) );
  HS65_LL_NOR4ABX2 U12280 ( .A(n10030), .B(n9982), .C(n9740), .D(n10186), .Z(
        n9741) );
  HS65_LL_NAND3X2 U12281 ( .A(n9743), .B(n9742), .C(n9741), .Z(n9744) );
  HS65_LL_MX41X4 U12282 ( .D0(n9747), .S0(n10221), .D1(n9746), .S1(n10308), 
        .D2(n9745), .S2(n10300), .D3(n9744), .S3(n10217), .Z(n9748) );
  HS65_LLS_XNOR2X3 U12283 ( .A(w0[2]), .B(n9748), .Z(n15024) );
  HS65_LL_MUX21I1X3 U12284 ( .D0(n15024), .D1(key[98]), .S0(n11617), .Z(
        \u0/N44 ) );
  HS65_LL_MUX21I1X3 U12285 ( .D0(n9749), .D1(key[109]), .S0(n15110), .Z(
        \u0/N55 ) );
  HS65_LL_NAND3X2 U12286 ( .A(n9752), .B(n9751), .C(n9750), .Z(n9753) );
  HS65_LL_NOR4ABX2 U12287 ( .A(n9755), .B(n9754), .C(n9879), .D(n9753), .Z(
        n10246) );
  HS65_LL_NAND4ABX3 U12288 ( .A(n9758), .B(n9757), .C(n10246), .D(n9756), .Z(
        n9788) );
  HS65_LL_NOR4ABX2 U12289 ( .A(n9761), .B(n9760), .C(n9759), .D(n9888), .Z(
        n9764) );
  HS65_LL_NOR4ABX2 U12290 ( .A(n9765), .B(n9764), .C(n9763), .D(n9762), .Z(
        n9785) );
  HS65_LL_NAND2X2 U12291 ( .A(n9910), .B(n9766), .Z(n10227) );
  HS65_LL_NOR4ABX2 U12292 ( .A(n9777), .B(n9768), .C(n9767), .D(n9900), .Z(
        n9769) );
  HS65_LL_NAND4ABX3 U12293 ( .A(n10249), .B(n10227), .C(n9770), .D(n9769), .Z(
        n9783) );
  HS65_LL_NOR4ABX2 U12294 ( .A(n9774), .B(n9773), .C(n9772), .D(n9771), .Z(
        n9781) );
  HS65_LL_OR2X4 U12295 ( .A(n9775), .B(n9880), .Z(n9776) );
  HS65_LL_NOR4ABX2 U12296 ( .A(n9778), .B(n9777), .C(n9776), .D(n9907), .Z(
        n9779) );
  HS65_LL_AOI13X2 U12297 ( .A(n9781), .B(n9780), .C(n9779), .D(n10257), .Z(
        n9782) );
  HS65_LL_CBI4I6X2 U12298 ( .A(n9906), .B(n9783), .C(n9919), .D(n9782), .Z(
        n9784) );
  HS65_LL_CBI4I1X3 U12299 ( .A(n9786), .B(n9785), .C(n10264), .D(n9784), .Z(
        n9787) );
  HS65_LL_AOI12X2 U12300 ( .A(n10260), .B(n9788), .C(n9787), .Z(n9789) );
  HS65_LLS_XOR2X3 U12301 ( .A(w0[22]), .B(n9789), .Z(n15028) );
  HS65_LL_MUX21I1X3 U12302 ( .D0(n15028), .D1(key[118]), .S0(n15783), .Z(
        \u0/N64 ) );
  HS65_LL_IVX2 U12303 ( .A(w0[10]), .Z(n15539) );
  HS65_LL_AOI112X2 U12304 ( .A(n9793), .B(n9792), .C(n9791), .D(n9790), .Z(
        n9796) );
  HS65_LL_NOR4ABX2 U12305 ( .A(n9797), .B(n9796), .C(n9795), .D(n9794), .Z(
        n9829) );
  HS65_LL_NAND3X2 U12306 ( .A(n9800), .B(n9799), .C(n9798), .Z(n9807) );
  HS65_LL_NOR4ABX2 U12307 ( .A(n9804), .B(n9803), .C(n9802), .D(n9801), .Z(
        n9805) );
  HS65_LL_NAND4ABX3 U12308 ( .A(n9808), .B(n9807), .C(n9806), .D(n9805), .Z(
        n9827) );
  HS65_LL_NOR4ABX2 U12309 ( .A(n9846), .B(n9811), .C(n9810), .D(n9809), .Z(
        n9824) );
  HS65_LL_NOR4ABX2 U12310 ( .A(n9824), .B(n9813), .C(n9833), .D(n9812), .Z(
        n9814) );
  HS65_LL_AOI13X2 U12311 ( .A(n9815), .B(n9814), .C(n9849), .D(n9866), .Z(
        n9826) );
  HS65_LL_NAND3X2 U12312 ( .A(n9860), .B(n9817), .C(n9816), .Z(n9818) );
  HS65_LL_NOR4ABX2 U12313 ( .A(n9821), .B(n9820), .C(n9819), .D(n9818), .Z(
        n9822) );
  HS65_LL_AOI13X2 U12314 ( .A(n9824), .B(n9823), .C(n9822), .D(n9854), .Z(
        n9825) );
  HS65_LL_AOI112X2 U12315 ( .A(n9873), .B(n9827), .C(n9826), .D(n9825), .Z(
        n9828) );
  HS65_LL_CBI4I1X3 U12316 ( .A(n9830), .B(n9829), .C(n9875), .D(n9828), .Z(
        n9831) );
  HS65_LL_MUXI21X2 U12317 ( .D0(w0[10]), .D1(n15539), .S0(n9831), .Z(n15034)
         );
  HS65_LL_MUX21I1X3 U12318 ( .D0(n15034), .D1(key[106]), .S0(n15110), .Z(
        \u0/N52 ) );
  HS65_LL_NAND2AX4 U12319 ( .A(n9833), .B(n9832), .Z(n9848) );
  HS65_LL_NAND4ABX3 U12320 ( .A(n9848), .B(n9836), .C(n9835), .D(n9834), .Z(
        n9837) );
  HS65_LL_NOR4ABX2 U12321 ( .A(n9840), .B(n9839), .C(n9838), .D(n9837), .Z(
        n9876) );
  HS65_LL_NOR4ABX2 U12322 ( .A(n9844), .B(n9843), .C(n9842), .D(n9841), .Z(
        n9845) );
  HS65_LL_NAND4ABX3 U12323 ( .A(n9848), .B(n9847), .C(n9846), .D(n9845), .Z(
        n9872) );
  HS65_LL_IVX2 U12324 ( .A(n9849), .Z(n9851) );
  HS65_LL_NOR4ABX2 U12325 ( .A(n9853), .B(n9852), .C(n9851), .D(n9850), .Z(
        n9855) );
  HS65_LL_AOI13X2 U12326 ( .A(n9857), .B(n9856), .C(n9855), .D(n9854), .Z(
        n9871) );
  HS65_LL_NOR4ABX2 U12327 ( .A(n9861), .B(n9860), .C(n9859), .D(n9858), .Z(
        n9865) );
  HS65_LL_NOR4ABX2 U12328 ( .A(n9865), .B(n9864), .C(n9863), .D(n9862), .Z(
        n9867) );
  HS65_LL_AOI13X2 U12329 ( .A(n9869), .B(n9868), .C(n9867), .D(n9866), .Z(
        n9870) );
  HS65_LL_AOI112X2 U12330 ( .A(n9873), .B(n9872), .C(n9871), .D(n9870), .Z(
        n9874) );
  HS65_LL_CBI4I1X3 U12331 ( .A(n9877), .B(n9876), .C(n9875), .D(n9874), .Z(
        n9878) );
  HS65_LLS_XNOR2X3 U12332 ( .A(w0[8]), .B(n9878), .Z(n15026) );
  HS65_LL_MUX21I1X3 U12333 ( .D0(n15026), .D1(key[104]), .S0(n15783), .Z(
        \u0/N50 ) );
  HS65_LL_IVX2 U12334 ( .A(w0[19]), .Z(n15257) );
  HS65_LL_NOR4ABX2 U12335 ( .A(n9882), .B(n9881), .C(n9880), .D(n9879), .Z(
        n9883) );
  HS65_LL_NAND4ABX3 U12336 ( .A(n9886), .B(n9885), .C(n9884), .D(n9883), .Z(
        n9921) );
  HS65_LL_AND2X4 U12337 ( .A(n9901), .B(n9887), .Z(n9893) );
  HS65_LL_NOR4ABX2 U12338 ( .A(n9891), .B(n9890), .C(n9889), .D(n9888), .Z(
        n9892) );
  HS65_LL_NAND4ABX3 U12339 ( .A(n10231), .B(n9894), .C(n9893), .D(n9892), .Z(
        n9897) );
  HS65_LL_NAND4ABX3 U12340 ( .A(n9898), .B(n9897), .C(n9896), .D(n9895), .Z(
        n9920) );
  HS65_LL_NOR4ABX2 U12341 ( .A(n9902), .B(n9901), .C(n9900), .D(n9899), .Z(
        n9903) );
  HS65_LL_NAND4ABX3 U12342 ( .A(n9906), .B(n9905), .C(n9904), .D(n9903), .Z(
        n9918) );
  HS65_LL_NOR4ABX2 U12343 ( .A(n9910), .B(n9909), .C(n9908), .D(n9907), .Z(
        n9911) );
  HS65_LL_NAND4ABX3 U12344 ( .A(n9914), .B(n9913), .C(n9912), .D(n9911), .Z(
        n9916) );
  HS65_LL_MX41X4 U12345 ( .D0(n9921), .S0(n10260), .D1(n9920), .S1(n9919), 
        .D2(n9918), .S2(n9917), .D3(n9916), .S3(n9915), .Z(n9922) );
  HS65_LL_MUXI21X2 U12346 ( .D0(w0[19]), .D1(n15257), .S0(n9922), .Z(n15037)
         );
  HS65_LL_MUX21I1X3 U12347 ( .D0(n15037), .D1(key[115]), .S0(n11617), .Z(
        \u0/N61 ) );
  HS65_LL_MUX21I1X3 U12348 ( .D0(n12148), .D1(n12148), .S0(w1[5]), .Z(N484) );
  HS65_LL_NOR4ABX2 U12349 ( .A(n9924), .B(n9923), .C(n9949), .D(n10019), .Z(
        n10286) );
  HS65_LL_NOR2X2 U12350 ( .A(n10270), .B(n9925), .Z(n10214) );
  HS65_LL_NAND3X2 U12351 ( .A(n10031), .B(n9926), .C(n10020), .Z(n10045) );
  HS65_LL_NOR4ABX2 U12352 ( .A(n10214), .B(n9927), .C(n10045), .D(n10201), .Z(
        n9928) );
  HS65_LL_NAND3X2 U12353 ( .A(n9929), .B(n10286), .C(n9928), .Z(n9956) );
  HS65_LL_NOR2X2 U12354 ( .A(n10213), .B(n10194), .Z(n10285) );
  HS65_LL_NAND4ABX3 U12355 ( .A(n9931), .B(n9930), .C(n10006), .D(n10285), .Z(
        n9932) );
  HS65_LL_NAND4ABX3 U12356 ( .A(n9933), .B(n9932), .C(n9979), .D(n9985), .Z(
        n9955) );
  HS65_LL_NOR2X2 U12357 ( .A(n9935), .B(n9934), .Z(n9964) );
  HS65_LL_NAND2X2 U12358 ( .A(n10020), .B(n10015), .Z(n10003) );
  HS65_LL_NOR3X1 U12359 ( .A(n10037), .B(n9973), .C(n10003), .Z(n9938) );
  HS65_LL_NOR4ABX2 U12360 ( .A(n9985), .B(n9938), .C(n9937), .D(n9936), .Z(
        n9939) );
  HS65_LL_NAND3X2 U12361 ( .A(n9964), .B(n9940), .C(n9939), .Z(n9954) );
  HS65_LL_CBI4I1X3 U12362 ( .A(n9944), .B(n9943), .C(n9942), .D(n9941), .Z(
        n9946) );
  HS65_LL_NAND4ABX3 U12363 ( .A(n9947), .B(n9946), .C(n10214), .D(n9945), .Z(
        n9952) );
  HS65_LL_NOR3X1 U12364 ( .A(n9950), .B(n9949), .C(n9948), .Z(n9971) );
  HS65_LL_NAND4ABX3 U12365 ( .A(n10209), .B(n9952), .C(n9971), .D(n9951), .Z(
        n9953) );
  HS65_LL_MX41X4 U12366 ( .D0(n9956), .S0(n10221), .D1(n9955), .S1(n10308), 
        .D2(n9954), .S2(n10300), .D3(n9953), .S3(n10217), .Z(n9957) );
  HS65_LLS_XNOR2X3 U12367 ( .A(w0[7]), .B(n9957), .Z(n15039) );
  HS65_LL_MUX21I1X3 U12368 ( .D0(n15039), .D1(key[103]), .S0(n11617), .Z(
        \u0/N49 ) );
  HS65_LL_IVX2 U12369 ( .A(w0[4]), .Z(n15438) );
  HS65_LL_NAND2X2 U12370 ( .A(n9958), .B(n10036), .Z(n10284) );
  HS65_LL_NOR2X2 U12371 ( .A(n10184), .B(n10284), .Z(n9992) );
  HS65_LL_IVX2 U12372 ( .A(n9986), .Z(n10296) );
  HS65_LL_NAND3X2 U12373 ( .A(n10296), .B(n9960), .C(n9959), .Z(n10289) );
  HS65_LL_NOR4ABX2 U12374 ( .A(n10182), .B(n9961), .C(n10270), .D(n10289), .Z(
        n9962) );
  HS65_LL_NAND4ABX3 U12375 ( .A(n10034), .B(n9963), .C(n9992), .D(n9962), .Z(
        n10000) );
  HS65_LL_NOR2X2 U12376 ( .A(n10290), .B(n10202), .Z(n9965) );
  HS65_LL_NAND4ABX3 U12377 ( .A(n9966), .B(n10284), .C(n9965), .D(n9964), .Z(
        n9967) );
  HS65_LL_NOR3X1 U12378 ( .A(n9968), .B(n10209), .C(n9967), .Z(n10306) );
  HS65_LL_NOR4ABX2 U12379 ( .A(n9969), .B(n10306), .C(n10292), .D(n10184), .Z(
        n10210) );
  HS65_LL_NAND2X2 U12380 ( .A(n9971), .B(n9970), .Z(n9993) );
  HS65_LL_NOR2X2 U12381 ( .A(n10196), .B(n9993), .Z(n10005) );
  HS65_LL_NOR4ABX2 U12382 ( .A(n10027), .B(n10199), .C(n10037), .D(n9972), .Z(
        n9975) );
  HS65_LL_NOR4ABX2 U12383 ( .A(n9976), .B(n9975), .C(n9974), .D(n9973), .Z(
        n9977) );
  HS65_LL_AOI13X2 U12384 ( .A(n10210), .B(n10005), .C(n9977), .D(n10295), .Z(
        n9999) );
  HS65_LL_NOR4ABX2 U12385 ( .A(n10197), .B(n9979), .C(n9993), .D(n9978), .Z(
        n9983) );
  HS65_LL_NOR4ABX2 U12386 ( .A(n9983), .B(n9982), .C(n9981), .D(n9980), .Z(
        n9997) );
  HS65_LL_NAND4ABX3 U12387 ( .A(n9986), .B(n10271), .C(n9985), .D(n9984), .Z(
        n9995) );
  HS65_LL_CB4I1X4 U12388 ( .A(n9990), .B(n9989), .C(n9988), .D(n9987), .Z(
        n9991) );
  HS65_LL_NAND4ABX3 U12389 ( .A(n9993), .B(n10209), .C(n9992), .D(n9991), .Z(
        n9994) );
  HS65_LL_OAI13X1 U12390 ( .A(n10029), .B(n9995), .C(n9994), .D(n10308), .Z(
        n9996) );
  HS65_LL_CBI4I1X3 U12391 ( .A(n10031), .B(n9997), .C(n10304), .D(n9996), .Z(
        n9998) );
  HS65_LL_AOI112X2 U12392 ( .A(n10300), .B(n10000), .C(n9999), .D(n9998), .Z(
        n10001) );
  HS65_LL_MUXI21X2 U12393 ( .D0(n15438), .D1(w0[4]), .S0(n10001), .Z(n15043)
         );
  HS65_LL_MUX21I1X3 U12394 ( .D0(n15043), .D1(key[100]), .S0(n15110), .Z(
        \u0/N46 ) );
  HS65_LL_NOR3AX2 U12395 ( .A(n10211), .B(n10003), .C(n10002), .Z(n10004) );
  HS65_LL_NAND3X2 U12396 ( .A(n10006), .B(n10005), .C(n10004), .Z(n10291) );
  HS65_LL_NAND4ABX3 U12397 ( .A(n10009), .B(n10284), .C(n10008), .D(n10007), 
        .Z(n10013) );
  HS65_LL_NAND2X2 U12398 ( .A(n10187), .B(n10010), .Z(n10012) );
  HS65_LL_NAND4ABX3 U12399 ( .A(n10014), .B(n10013), .C(n10012), .D(n10011), 
        .Z(n10025) );
  HS65_LL_NAND2X2 U12400 ( .A(n10016), .B(n10015), .Z(n10277) );
  HS65_LL_NOR4ABX2 U12401 ( .A(n10018), .B(n10017), .C(n10272), .D(n10277), 
        .Z(n10021) );
  HS65_LL_NOR4ABX2 U12402 ( .A(n10021), .B(n10020), .C(n10184), .D(n10019), 
        .Z(n10022) );
  HS65_LL_AOI13X2 U12403 ( .A(n10027), .B(n10023), .C(n10022), .D(n10304), .Z(
        n10024) );
  HS65_LL_CBI4I6X2 U12404 ( .A(n10291), .B(n10025), .C(n10300), .D(n10024), 
        .Z(n10049) );
  HS65_LL_NAND4ABX3 U12405 ( .A(n10029), .B(n10028), .C(n10027), .D(n10026), 
        .Z(n10035) );
  HS65_LL_NAND4ABX3 U12406 ( .A(n10194), .B(n10032), .C(n10031), .D(n10030), 
        .Z(n10033) );
  HS65_LL_OAI13X1 U12407 ( .A(n10035), .B(n10034), .C(n10033), .D(n10217), .Z(
        n10048) );
  HS65_LL_NAND2AX4 U12408 ( .A(n10037), .B(n10036), .Z(n10193) );
  HS65_LL_NAND3X2 U12409 ( .A(n10040), .B(n10039), .C(n10038), .Z(n10043) );
  HS65_LL_NAND4ABX3 U12410 ( .A(n10193), .B(n10043), .C(n10042), .D(n10041), 
        .Z(n10044) );
  HS65_LL_OAI13X1 U12411 ( .A(n10046), .B(n10045), .C(n10044), .D(n10308), .Z(
        n10047) );
  HS65_LL_NAND3X2 U12412 ( .A(n10049), .B(n10048), .C(n10047), .Z(n10050) );
  HS65_LLS_XNOR2X3 U12413 ( .A(w0[0]), .B(n10050), .Z(n15041) );
  HS65_LL_MUX21I1X3 U12414 ( .D0(n15041), .D1(key[96]), .S0(n11617), .Z(
        \u0/N42 ) );
  HS65_LL_NOR2X2 U12415 ( .A(n11025), .B(n10056), .Z(n13370) );
  HS65_LL_NOR2X2 U12416 ( .A(n10960), .B(n10051), .Z(n11051) );
  HS65_LL_NOR3X1 U12417 ( .A(n11060), .B(n13370), .C(n11051), .Z(n10730) );
  HS65_LL_NAND2X2 U12418 ( .A(n10052), .B(n10612), .Z(n10738) );
  HS65_LL_NOR4ABX2 U12419 ( .A(n10738), .B(n13397), .C(n10054), .D(n10053), 
        .Z(n10055) );
  HS65_LL_NAND3X2 U12420 ( .A(n10730), .B(n10069), .C(n10055), .Z(n13396) );
  HS65_LL_NAND2X2 U12421 ( .A(n10626), .B(n11042), .Z(n10643) );
  HS65_LL_NOR2X2 U12422 ( .A(n10056), .B(n10958), .Z(n11044) );
  HS65_LL_IVX2 U12423 ( .A(n11045), .Z(n13387) );
  HS65_LL_NOR2X2 U12424 ( .A(n10736), .B(n13387), .Z(n13372) );
  HS65_LL_NAND4ABX3 U12425 ( .A(n11044), .B(n10073), .C(n13372), .D(n13367), 
        .Z(n10057) );
  HS65_LL_NOR3X1 U12426 ( .A(n10716), .B(n10729), .C(n10057), .Z(n10820) );
  HS65_LL_NAND4ABX3 U12427 ( .A(n10951), .B(n10643), .C(n10820), .D(n10948), 
        .Z(n10058) );
  HS65_LL_NOR2X2 U12428 ( .A(n10811), .B(n10955), .Z(n10064) );
  HS65_LL_NOR3AX2 U12429 ( .A(n10064), .B(n11064), .C(n10829), .Z(n11034) );
  HS65_LL_NAND2X2 U12430 ( .A(sa12[5]), .B(n10954), .Z(n10732) );
  HS65_LL_NAND4ABX3 U12431 ( .A(n10934), .B(n10058), .C(n11034), .D(n10732), 
        .Z(n10083) );
  HS65_LL_NOR2X2 U12432 ( .A(n11060), .B(n10606), .Z(n11023) );
  HS65_LL_NOR2X2 U12433 ( .A(n10743), .B(n10070), .Z(n10621) );
  HS65_LL_NOR2X2 U12434 ( .A(n13400), .B(n10716), .Z(n13381) );
  HS65_LL_NOR2X2 U12435 ( .A(n10711), .B(n11051), .Z(n10834) );
  HS65_LL_NAND4ABX3 U12436 ( .A(n10934), .B(n13383), .C(n10807), .D(n10834), 
        .Z(n10059) );
  HS65_LL_NOR4ABX2 U12437 ( .A(n10621), .B(n13381), .C(n10643), .D(n10059), 
        .Z(n11062) );
  HS65_LL_NOR4ABX2 U12438 ( .A(n11023), .B(n11062), .C(n10620), .D(n10073), 
        .Z(n10081) );
  HS65_LL_NOR2X2 U12439 ( .A(n10060), .B(n10958), .Z(n10062) );
  HS65_LL_NOR3X1 U12440 ( .A(n10962), .B(n10062), .C(n10061), .Z(n11056) );
  HS65_LL_AND2X4 U12441 ( .A(n10742), .B(n10826), .Z(n10728) );
  HS65_LL_NOR2X2 U12442 ( .A(n10960), .B(n10629), .Z(n13388) );
  HS65_LL_NOR4ABX2 U12443 ( .A(n10738), .B(n10728), .C(n11033), .D(n13388), 
        .Z(n10063) );
  HS65_LL_NAND3X2 U12444 ( .A(n10064), .B(n11035), .C(n10063), .Z(n10759) );
  HS65_LL_NAND4ABX3 U12445 ( .A(n11048), .B(n10759), .C(n10065), .D(n11057), 
        .Z(n10066) );
  HS65_LL_NOR4ABX2 U12446 ( .A(n11056), .B(n13397), .C(n10931), .D(n10066), 
        .Z(n10080) );
  HS65_LL_IVX2 U12447 ( .A(n10081), .Z(n10078) );
  HS65_LL_NAND2X2 U12448 ( .A(n10617), .B(n11030), .Z(n10950) );
  HS65_LL_NOR2X2 U12449 ( .A(n13370), .B(n11048), .Z(n10640) );
  HS65_LL_NAND4ABX3 U12450 ( .A(n10931), .B(n10825), .C(n10640), .D(n11022), 
        .Z(n10067) );
  HS65_LL_NOR2X2 U12451 ( .A(n11043), .B(n11064), .Z(n10712) );
  HS65_LL_NAND4ABX3 U12452 ( .A(n13388), .B(n10067), .C(n10712), .D(n10826), 
        .Z(n13378) );
  HS65_LL_NOR4ABX2 U12453 ( .A(n10725), .B(n11052), .C(n13365), .D(n13386), 
        .Z(n10068) );
  HS65_LL_NAND4ABX3 U12454 ( .A(n10950), .B(n13378), .C(n10069), .D(n10068), 
        .Z(n10077) );
  HS65_LL_IVX2 U12455 ( .A(n11044), .Z(n10717) );
  HS65_LL_NOR4ABX2 U12456 ( .A(n10717), .B(n10725), .C(n10619), .D(n10070), 
        .Z(n11031) );
  HS65_LL_NOR3AX2 U12457 ( .A(n10948), .B(n10833), .C(n13388), .Z(n11049) );
  HS65_LL_NOR3X1 U12458 ( .A(n13365), .B(n10955), .C(n10624), .Z(n10074) );
  HS65_LL_NOR4ABX2 U12459 ( .A(n10071), .B(n11042), .C(n10620), .D(n10825), 
        .Z(n10072) );
  HS65_LL_NAND3X2 U12460 ( .A(n13368), .B(n11056), .C(n10072), .Z(n10754) );
  HS65_LL_NOR4ABX2 U12461 ( .A(n10074), .B(n10807), .C(n10073), .D(n10754), 
        .Z(n10075) );
  HS65_LL_AOI13X2 U12462 ( .A(n11031), .B(n11049), .C(n10075), .D(n10756), .Z(
        n10076) );
  HS65_LL_CBI4I6X2 U12463 ( .A(n10078), .B(n10077), .C(n11068), .D(n10076), 
        .Z(n10079) );
  HS65_LL_CBI4I1X3 U12464 ( .A(n10081), .B(n10080), .C(n10750), .D(n10079), 
        .Z(n10082) );
  HS65_LL_CBI4I6X2 U12465 ( .A(n13396), .B(n10083), .C(n13401), .D(n10082), 
        .Z(n14647) );
  HS65_LL_MUX21I1X3 U12466 ( .D0(n14647), .D1(n14647), .S0(w1[18]), .Z(N423)
         );
  HS65_LL_MUX21I1X3 U12467 ( .D0(n10084), .D1(key[121]), .S0(n15110), .Z(
        \u0/N67 ) );
  HS65_LLS_XNOR2X3 U12468 ( .A(w1[18]), .B(n10085), .Z(n15827) );
  HS65_LLS_XNOR2X3 U12469 ( .A(w2[18]), .B(n15827), .Z(n15784) );
  HS65_LL_MUX21I1X3 U12470 ( .D0(n15784), .D1(key[50]), .S0(n15110), .Z(
        \u0/N192 ) );
  HS65_LL_MUX21I1X3 U12471 ( .D0(n10086), .D1(key[77]), .S0(n11617), .Z(
        \u0/N121 ) );
  HS65_LL_AOI12X2 U12472 ( .A(n12922), .B(n10131), .C(n12453), .Z(n11319) );
  HS65_LL_IVX2 U12473 ( .A(n10120), .Z(n12476) );
  HS65_LL_IVX2 U12474 ( .A(n11761), .Z(n12489) );
  HS65_LL_NAND2X2 U12475 ( .A(n10087), .B(n11340), .Z(n10115) );
  HS65_LL_NAND2X2 U12476 ( .A(n12489), .B(n10115), .Z(n11330) );
  HS65_LL_AOI112X2 U12477 ( .A(n11309), .B(n10088), .C(n12476), .D(n11330), 
        .Z(n10089) );
  HS65_LL_NAND4ABX3 U12478 ( .A(n11334), .B(n11335), .C(n11319), .D(n10089), 
        .Z(n12934) );
  HS65_LL_NAND2AX4 U12479 ( .A(n12504), .B(n10090), .Z(n11670) );
  HS65_LL_NOR2X2 U12480 ( .A(n10117), .B(n10091), .Z(n11756) );
  HS65_LL_AOI12X2 U12481 ( .A(n10130), .B(n12930), .C(n12441), .Z(n11763) );
  HS65_LL_NOR2X2 U12482 ( .A(n10112), .B(n10091), .Z(n11738) );
  HS65_LL_NOR3X1 U12483 ( .A(n11744), .B(n12462), .C(n11738), .Z(n11316) );
  HS65_LL_NAND4ABX3 U12484 ( .A(n12469), .B(n11756), .C(n11763), .D(n11316), 
        .Z(n10094) );
  HS65_LL_NAND2X2 U12485 ( .A(n11665), .B(n11739), .Z(n12438) );
  HS65_LL_NOR3X1 U12486 ( .A(n12936), .B(n10092), .C(n12438), .Z(n10106) );
  HS65_LL_NAND2AX4 U12487 ( .A(n10098), .B(n10123), .Z(n12935) );
  HS65_LL_NOR2AX3 U12488 ( .A(n12448), .B(n12935), .Z(n10105) );
  HS65_LL_NAND2X2 U12489 ( .A(n10105), .B(n11313), .Z(n11333) );
  HS65_LL_NOR2X2 U12490 ( .A(n10093), .B(n11333), .Z(n11678) );
  HS65_LL_NAND4ABX3 U12491 ( .A(n11670), .B(n10094), .C(n10106), .D(n11678), 
        .Z(n10142) );
  HS65_LL_IVX2 U12492 ( .A(n12947), .Z(n12540) );
  HS65_LL_NOR4ABX2 U12493 ( .A(n12473), .B(n11313), .C(n11747), .D(n10095), 
        .Z(n12909) );
  HS65_LL_NAND4ABX3 U12494 ( .A(n10096), .B(n12462), .C(n12477), .D(n12515), 
        .Z(n10097) );
  HS65_LL_NOR3X1 U12495 ( .A(n10098), .B(n12460), .C(n10097), .Z(n11741) );
  HS65_LL_NOR2X2 U12496 ( .A(n10099), .B(n12498), .Z(n12454) );
  HS65_LL_NAND2X2 U12497 ( .A(n11311), .B(n11309), .Z(n12470) );
  HS65_LL_OAI112X1 U12498 ( .A(n10101), .B(n10100), .C(n12454), .D(n12470), 
        .Z(n10102) );
  HS65_LL_NOR2X2 U12499 ( .A(n11743), .B(n10127), .Z(n11683) );
  HS65_LL_NAND4ABX3 U12500 ( .A(n11318), .B(n10102), .C(n12911), .D(n11683), 
        .Z(n10103) );
  HS65_LL_NOR4ABX2 U12501 ( .A(n12909), .B(n11741), .C(n10104), .D(n10103), 
        .Z(n10140) );
  HS65_LL_NAND2X2 U12502 ( .A(n10106), .B(n10105), .Z(n12519) );
  HS65_LL_OAI21X2 U12503 ( .A(n10108), .B(n11340), .C(n10107), .Z(n12466) );
  HS65_LL_NAND3X2 U12504 ( .A(n10109), .B(n11683), .C(n12466), .Z(n10113) );
  HS65_LL_NOR2X2 U12505 ( .A(n10111), .B(n10110), .Z(n12937) );
  HS65_LL_NOR2X2 U12506 ( .A(n10112), .B(n10133), .Z(n12503) );
  HS65_LL_NAND2AX4 U12507 ( .A(n12503), .B(n10115), .Z(n12439) );
  HS65_LL_NOR2X2 U12508 ( .A(n12937), .B(n12439), .Z(n11672) );
  HS65_LL_NAND4ABX3 U12509 ( .A(n12535), .B(n10113), .C(n12509), .D(n11672), 
        .Z(n10114) );
  HS65_LL_OAI21X2 U12510 ( .A(n12519), .B(n10114), .C(n12945), .Z(n10139) );
  HS65_LL_NAND2AX4 U12511 ( .A(n12505), .B(n10115), .Z(n12907) );
  HS65_LL_NAND2X2 U12512 ( .A(n11661), .B(n10116), .Z(n11328) );
  HS65_LL_NOR2X2 U12513 ( .A(n10118), .B(n10117), .Z(n11688) );
  HS65_LL_NAND2X2 U12514 ( .A(sa22[1]), .B(n11688), .Z(n12516) );
  HS65_LL_OAI21X2 U12515 ( .A(n11675), .B(n10119), .C(n12516), .Z(n12468) );
  HS65_LL_NAND3X2 U12516 ( .A(sa22[6]), .B(n11309), .C(n11667), .Z(n12919) );
  HS65_LL_NAND2X2 U12517 ( .A(n10120), .B(n12919), .Z(n11755) );
  HS65_LL_NOR2AX3 U12518 ( .A(n10121), .B(n11310), .Z(n11690) );
  HS65_LL_NAND3AX3 U12519 ( .A(n11756), .B(n11690), .C(n10122), .Z(n12529) );
  HS65_LL_NOR4ABX2 U12520 ( .A(n12911), .B(n10123), .C(n11755), .D(n12529), 
        .Z(n10136) );
  HS65_LL_NOR2X2 U12521 ( .A(n11323), .B(n10124), .Z(n11736) );
  HS65_LL_IVX2 U12522 ( .A(n11747), .Z(n12531) );
  HS65_LL_NAND3X2 U12523 ( .A(n10125), .B(n12470), .C(n12531), .Z(n10126) );
  HS65_LL_NOR3X1 U12524 ( .A(n10127), .B(n11736), .C(n10126), .Z(n12442) );
  HS65_LL_NOR2X2 U12525 ( .A(n10129), .B(n10128), .Z(n12499) );
  HS65_LL_NAND2X2 U12526 ( .A(n11680), .B(n12477), .Z(n12916) );
  HS65_LL_CBI4I6X2 U12527 ( .A(n10131), .B(n12499), .C(n10130), .D(n12916), 
        .Z(n10132) );
  HS65_LL_OAI112X1 U12528 ( .A(n10134), .B(n10133), .C(n12442), .D(n10132), 
        .Z(n12926) );
  HS65_LL_NOR4ABX2 U12529 ( .A(n10136), .B(n12501), .C(n10135), .D(n12926), 
        .Z(n11342) );
  HS65_LL_NOR4X4 U12530 ( .A(n11738), .B(n12441), .C(n11743), .D(n12498), .Z(
        n12494) );
  HS65_LL_NAND4ABX3 U12531 ( .A(n11328), .B(n12468), .C(n11342), .D(n12494), 
        .Z(n10137) );
  HS65_LL_OAI13X1 U12532 ( .A(n11308), .B(n12907), .C(n10137), .D(n12951), .Z(
        n10138) );
  HS65_LL_OAI112X1 U12533 ( .A(n10140), .B(n11339), .C(n10139), .D(n10138), 
        .Z(n10141) );
  HS65_LL_CBI4I6X2 U12534 ( .A(n12934), .B(n10142), .C(n12540), .D(n10141), 
        .Z(n14633) );
  HS65_LL_MUX21I1X3 U12535 ( .D0(n14633), .D1(n14633), .S0(w0[8]), .Z(N449) );
  HS65_LL_NAND2X2 U12536 ( .A(n10153), .B(n12169), .Z(n12833) );
  HS65_LL_NOR2X2 U12537 ( .A(n10885), .B(n11129), .Z(n12818) );
  HS65_LL_NAND2X2 U12538 ( .A(n10164), .B(n10143), .Z(n12163) );
  HS65_LL_NOR4ABX2 U12539 ( .A(n10144), .B(n12163), .C(n14655), .D(n14649), 
        .Z(n10148) );
  HS65_LL_NOR2X2 U12540 ( .A(n10146), .B(n10145), .Z(n12181) );
  HS65_LL_NAND2X2 U12541 ( .A(n10909), .B(n10889), .Z(n10919) );
  HS65_LL_NOR4ABX2 U12542 ( .A(n10148), .B(n10147), .C(n12181), .D(n10919), 
        .Z(n14689) );
  HS65_LL_NAND4ABX3 U12543 ( .A(n10149), .B(n12180), .C(n12818), .D(n14689), 
        .Z(n10150) );
  HS65_LL_NAND4ABX3 U12544 ( .A(n12833), .B(n10150), .C(n12178), .D(n12827), 
        .Z(n10181) );
  HS65_LL_NAND3X2 U12545 ( .A(n14651), .B(n10917), .C(n10906), .Z(n10151) );
  HS65_LL_NOR3X1 U12546 ( .A(n12819), .B(n10152), .C(n10151), .Z(n11135) );
  HS65_LL_IVX2 U12547 ( .A(n10153), .Z(n10911) );
  HS65_LL_NOR2X2 U12548 ( .A(n10911), .B(n10154), .Z(n12164) );
  HS65_LL_NOR2X2 U12549 ( .A(n10155), .B(n10171), .Z(n14657) );
  HS65_LL_NAND3AX3 U12550 ( .A(n14657), .B(n10157), .C(n10156), .Z(n12183) );
  HS65_LL_AOI112X2 U12551 ( .A(n10159), .B(n10158), .C(n14655), .D(n12183), 
        .Z(n10162) );
  HS65_LL_NAND2AX4 U12552 ( .A(n10168), .B(n12184), .Z(n10160) );
  HS65_LL_NOR4ABX2 U12553 ( .A(n12164), .B(n10162), .C(n10161), .D(n10160), 
        .Z(n10179) );
  HS65_LL_NOR2X2 U12554 ( .A(n14655), .B(n12813), .Z(n12828) );
  HS65_LL_NAND2X2 U12555 ( .A(n12178), .B(n12830), .Z(n11123) );
  HS65_LL_AOI13X2 U12556 ( .A(sa30[5]), .B(n10164), .C(n10163), .D(n11123), 
        .Z(n10166) );
  HS65_LL_NAND2X2 U12557 ( .A(n12177), .B(n10901), .Z(n11140) );
  HS65_LL_NOR4ABX2 U12558 ( .A(n14667), .B(n10166), .C(n10165), .D(n11140), 
        .Z(n12816) );
  HS65_LL_NAND4ABX3 U12559 ( .A(n10168), .B(n10167), .C(n12816), .D(n12184), 
        .Z(n10175) );
  HS65_LL_NOR4ABX2 U12560 ( .A(n12851), .B(n10916), .C(n10175), .D(n10169), 
        .Z(n10170) );
  HS65_LL_NAND3X2 U12561 ( .A(n12828), .B(n14673), .C(n10170), .Z(n10177) );
  HS65_LL_NOR2X2 U12562 ( .A(n10908), .B(n10171), .Z(n11130) );
  HS65_LL_NOR2X2 U12563 ( .A(n10900), .B(n11130), .Z(n12836) );
  HS65_LL_NAND2X2 U12564 ( .A(n12821), .B(n12850), .Z(n14669) );
  HS65_LL_NOR4ABX2 U12565 ( .A(n12836), .B(n11118), .C(n11125), .D(n14669), 
        .Z(n10172) );
  HS65_LL_NAND3X2 U12566 ( .A(n10172), .B(n10923), .C(n12174), .Z(n11137) );
  HS65_LL_NOR2X2 U12567 ( .A(n12834), .B(n12819), .Z(n12858) );
  HS65_LL_NOR4ABX2 U12568 ( .A(n10173), .B(n10909), .C(n12156), .D(n12176), 
        .Z(n10174) );
  HS65_LL_NAND4ABX3 U12569 ( .A(n10175), .B(n11137), .C(n12858), .D(n10174), 
        .Z(n10176) );
  HS65_LL_AOI22X1 U12570 ( .A(n14685), .B(n10177), .C(n14691), .D(n10176), .Z(
        n10178) );
  HS65_LL_CBI4I1X3 U12571 ( .A(n11135), .B(n10179), .C(n14687), .D(n10178), 
        .Z(n10180) );
  HS65_LL_CBI4I6X2 U12572 ( .A(n10886), .B(n10181), .C(n14683), .D(n10180), 
        .Z(n14854) );
  HS65_LL_MUX21I1X3 U12573 ( .D0(n14854), .D1(n14854), .S0(w1[2]), .Z(N487) );
  HS65_LL_IVX2 U12574 ( .A(w0[3]), .Z(n15440) );
  HS65_LL_NAND4ABX3 U12575 ( .A(n10273), .B(n10184), .C(n10183), .D(n10182), 
        .Z(n10185) );
  HS65_LL_AOI112X2 U12576 ( .A(n10188), .B(n10187), .C(n10186), .D(n10185), 
        .Z(n10189) );
  HS65_LL_NAND3X2 U12577 ( .A(n10274), .B(n10190), .C(n10189), .Z(n10222) );
  HS65_LL_NAND4ABX3 U12578 ( .A(n10194), .B(n10193), .C(n10192), .D(n10191), 
        .Z(n10195) );
  HS65_LL_NOR4ABX2 U12579 ( .A(n10198), .B(n10197), .C(n10196), .D(n10195), 
        .Z(n10200) );
  HS65_LL_NAND4ABX3 U12580 ( .A(n10202), .B(n10201), .C(n10200), .D(n10199), 
        .Z(n10220) );
  HS65_LL_NOR4ABX2 U12581 ( .A(n10206), .B(n10205), .C(n10204), .D(n10203), 
        .Z(n10207) );
  HS65_LL_NAND4ABX3 U12582 ( .A(n10302), .B(n10209), .C(n10208), .D(n10207), 
        .Z(n10219) );
  HS65_LL_NAND4ABX3 U12583 ( .A(n10213), .B(n10212), .C(n10211), .D(n10210), 
        .Z(n10215) );
  HS65_LL_NAND4ABX3 U12584 ( .A(n10216), .B(n10215), .C(n10288), .D(n10214), 
        .Z(n10218) );
  HS65_LL_MX41X4 U12585 ( .D0(n10222), .S0(n10221), .D1(n10220), .S1(n10308), 
        .D2(n10219), .S2(n10300), .D3(n10218), .S3(n10217), .Z(n10223) );
  HS65_LL_MUXI21X2 U12586 ( .D0(w0[3]), .D1(n15440), .S0(n10223), .Z(n15093)
         );
  HS65_LL_MUX21I1X3 U12587 ( .D0(n15093), .D1(key[99]), .S0(n15783), .Z(
        \u0/N45 ) );
  HS65_LL_NOR4ABX2 U12588 ( .A(n10233), .B(n10226), .C(n10225), .D(n10224), 
        .Z(n10228) );
  HS65_LL_NOR4ABX2 U12589 ( .A(n10229), .B(n10228), .C(n10236), .D(n10227), 
        .Z(n10265) );
  HS65_LL_NOR4ABX2 U12590 ( .A(n10233), .B(n10232), .C(n10231), .D(n10230), 
        .Z(n10234) );
  HS65_LL_NAND4ABX3 U12591 ( .A(n10237), .B(n10236), .C(n10235), .D(n10234), 
        .Z(n10261) );
  HS65_LL_NOR2X2 U12592 ( .A(w3[9]), .B(n10238), .Z(n10241) );
  HS65_LL_NAND4ABX3 U12593 ( .A(n10242), .B(n10241), .C(n10240), .D(n10239), 
        .Z(n10243) );
  HS65_LL_NOR4ABX2 U12594 ( .A(n10246), .B(n10245), .C(n10244), .D(n10243), 
        .Z(n10258) );
  HS65_LL_NAND4ABX3 U12595 ( .A(n10250), .B(n10249), .C(n10248), .D(n10247), 
        .Z(n10251) );
  HS65_LL_NOR4ABX2 U12596 ( .A(n10254), .B(n10253), .C(n10252), .D(n10251), 
        .Z(n10256) );
  HS65_LL_OAI22X1 U12597 ( .A(n10258), .B(n10257), .C(n10256), .D(n10255), .Z(
        n10259) );
  HS65_LL_CBI4I6X2 U12598 ( .A(n10262), .B(n10261), .C(n10260), .D(n10259), 
        .Z(n10263) );
  HS65_LL_CBI4I1X3 U12599 ( .A(n10266), .B(n10265), .C(n10264), .D(n10263), 
        .Z(n10267) );
  HS65_LLS_XNOR2X3 U12600 ( .A(w0[16]), .B(n10267), .Z(n15095) );
  HS65_LL_MUX21I1X3 U12601 ( .D0(n15095), .D1(key[112]), .S0(n15110), .Z(
        \u0/N58 ) );
  HS65_LL_NAND4ABX3 U12602 ( .A(n10271), .B(n10270), .C(n10269), .D(n10268), 
        .Z(n10276) );
  HS65_LL_NOR2X2 U12603 ( .A(n10273), .B(n10272), .Z(n10275) );
  HS65_LL_NAND4ABX3 U12604 ( .A(n10277), .B(n10276), .C(n10275), .D(n10274), 
        .Z(n10309) );
  HS65_LL_NAND3X2 U12605 ( .A(n10279), .B(n10278), .C(n10293), .Z(n10280) );
  HS65_LL_NOR4ABX2 U12606 ( .A(n10283), .B(n10282), .C(n10281), .D(n10280), 
        .Z(n10305) );
  HS65_LL_NOR4ABX2 U12607 ( .A(n10286), .B(n10285), .C(n10284), .D(n10310), 
        .Z(n10287) );
  HS65_LL_NAND4ABX3 U12608 ( .A(n10290), .B(n10289), .C(n10288), .D(n10287), 
        .Z(n10301) );
  HS65_LL_NOR4ABX2 U12609 ( .A(n10294), .B(n10293), .C(n10292), .D(n10291), 
        .Z(n10298) );
  HS65_LL_AOI13X2 U12610 ( .A(n10298), .B(n10297), .C(n10296), .D(n10295), .Z(
        n10299) );
  HS65_LL_CBI4I6X2 U12611 ( .A(n10302), .B(n10301), .C(n10300), .D(n10299), 
        .Z(n10303) );
  HS65_LL_CBI4I1X3 U12612 ( .A(n10306), .B(n10305), .C(n10304), .D(n10303), 
        .Z(n10307) );
  HS65_LL_CBI4I6X2 U12613 ( .A(n10310), .B(n10309), .C(n10308), .D(n10307), 
        .Z(n10311) );
  HS65_LLS_XOR2X3 U12614 ( .A(w0[6]), .B(n10311), .Z(n15097) );
  HS65_LL_MUX21I1X3 U12615 ( .D0(n15097), .D1(key[102]), .S0(n15110), .Z(
        \u0/N48 ) );
  HS65_LL_NOR2X2 U12616 ( .A(n10312), .B(n10469), .Z(n15079) );
  HS65_LL_NOR2X2 U12617 ( .A(n10410), .B(n10347), .Z(n10513) );
  HS65_LL_NOR2X2 U12618 ( .A(n10373), .B(n15077), .Z(n10465) );
  HS65_LL_NOR4ABX2 U12619 ( .A(n10465), .B(n10446), .C(n10370), .D(n10313), 
        .Z(n10314) );
  HS65_LL_NAND3X2 U12620 ( .A(n15079), .B(n10513), .C(n10314), .Z(n10501) );
  HS65_LL_IVX2 U12621 ( .A(n10332), .Z(n10508) );
  HS65_LL_NAND2X2 U12622 ( .A(n10508), .B(n10450), .Z(n10420) );
  HS65_LL_IVX2 U12623 ( .A(n10420), .Z(n10328) );
  HS65_LL_NAND4ABX3 U12624 ( .A(n10316), .B(n10382), .C(n10328), .D(n10315), 
        .Z(n10389) );
  HS65_LL_NOR4ABX2 U12625 ( .A(n10317), .B(n10494), .C(n15068), .D(n10336), 
        .Z(n10318) );
  HS65_LL_NAND4ABX3 U12626 ( .A(n10501), .B(n10389), .C(n10319), .D(n10318), 
        .Z(n10357) );
  HS65_LL_NOR2X2 U12627 ( .A(n10340), .B(n10320), .Z(n10458) );
  HS65_LL_NOR2X2 U12628 ( .A(n10456), .B(n10495), .Z(n10348) );
  HS65_LL_IVX2 U12629 ( .A(n10486), .Z(n15057) );
  HS65_LL_NOR4ABX2 U12630 ( .A(n10458), .B(n10348), .C(n10485), .D(n15057), 
        .Z(n10330) );
  HS65_LL_NOR2X2 U12631 ( .A(n10382), .B(n10321), .Z(n10512) );
  HS65_LL_IVX2 U12632 ( .A(n10322), .Z(n10325) );
  HS65_LL_NAND2X2 U12633 ( .A(n10323), .B(n10455), .Z(n15076) );
  HS65_LL_AOI112X2 U12634 ( .A(n10325), .B(n10324), .C(n10406), .D(n15076), 
        .Z(n10327) );
  HS65_LL_IVX2 U12635 ( .A(n10346), .Z(n15050) );
  HS65_LL_NOR3X1 U12636 ( .A(n10417), .B(n10326), .C(n10484), .Z(n15052) );
  HS65_LL_IVX2 U12637 ( .A(n10453), .Z(n10528) );
  HS65_LL_NAND2X2 U12638 ( .A(n15052), .B(n10528), .Z(n10339) );
  HS65_LL_NOR4ABX2 U12639 ( .A(n10328), .B(n10327), .C(n15050), .D(n10339), 
        .Z(n10329) );
  HS65_LL_AOI13X2 U12640 ( .A(n10330), .B(n10512), .C(n10329), .D(n10535), .Z(
        n10356) );
  HS65_LL_NOR2X2 U12641 ( .A(n10409), .B(n10331), .Z(n15063) );
  HS65_LL_NOR2X2 U12642 ( .A(n10511), .B(n10332), .Z(n10337) );
  HS65_LL_NOR2AX3 U12643 ( .A(n10412), .B(n10382), .Z(n15078) );
  HS65_LL_NAND4ABX3 U12644 ( .A(n10339), .B(n10334), .C(n10333), .D(n15078), 
        .Z(n10335) );
  HS65_LL_NOR4ABX2 U12645 ( .A(n10465), .B(n10337), .C(n10336), .D(n10335), 
        .Z(n10354) );
  HS65_LL_NOR2X2 U12646 ( .A(n15058), .B(n15068), .Z(n10530) );
  HS65_LL_NAND3X2 U12647 ( .A(n10338), .B(n10530), .C(n10446), .Z(n10351) );
  HS65_LL_IVX2 U12648 ( .A(n10370), .Z(n10411) );
  HS65_LL_NAND2X2 U12649 ( .A(n10362), .B(n10411), .Z(n10463) );
  HS65_LL_NOR2X2 U12650 ( .A(n10464), .B(n10339), .Z(n10379) );
  HS65_LL_NOR4ABX2 U12651 ( .A(n10342), .B(n10341), .C(n10340), .D(n15062), 
        .Z(n10413) );
  HS65_LL_NOR4ABX2 U12652 ( .A(n10344), .B(n10413), .C(n10343), .D(n10420), 
        .Z(n10345) );
  HS65_LL_IVX2 U12653 ( .A(n10449), .Z(n10387) );
  HS65_LL_NAND3X2 U12654 ( .A(n10346), .B(n10345), .C(n10387), .Z(n10369) );
  HS65_LL_NOR4ABX2 U12655 ( .A(n10349), .B(n10348), .C(n10347), .D(n10369), 
        .Z(n10470) );
  HS65_LL_NAND4ABX3 U12656 ( .A(n10502), .B(n10463), .C(n10379), .D(n10470), 
        .Z(n10350) );
  HS65_LL_OAI13X1 U12657 ( .A(n10352), .B(n10351), .C(n10350), .D(n15088), .Z(
        n10353) );
  HS65_LL_CBI4I1X3 U12658 ( .A(n15063), .B(n10354), .C(n10527), .D(n10353), 
        .Z(n10355) );
  HS65_LL_AOI112X2 U12659 ( .A(n15084), .B(n10357), .C(n10356), .D(n10355), 
        .Z(n10358) );
  HS65_LLS_XOR3X2 U12660 ( .A(n10358), .B(\u0/rcon [28]), .C(w0[28]), .Z(
        n15099) );
  HS65_LL_MUX21I1X3 U12661 ( .D0(n15099), .D1(key[124]), .S0(n11617), .Z(
        \u0/N70 ) );
  HS65_LL_MUX21I1X3 U12662 ( .D0(n10359), .D1(key[125]), .S0(n15110), .Z(
        \u0/N71 ) );
  HS65_LL_NAND4ABX3 U12663 ( .A(n10415), .B(n10360), .C(n10478), .D(n10516), 
        .Z(n10401) );
  HS65_LL_NOR3X1 U12664 ( .A(n10453), .B(n15058), .C(n15057), .Z(n10427) );
  HS65_LL_NAND2X2 U12665 ( .A(n10522), .B(n15051), .Z(n10408) );
  HS65_LL_NAND3X2 U12666 ( .A(n10362), .B(n10361), .C(n10381), .Z(n10505) );
  HS65_LL_NOR3AX2 U12667 ( .A(n10363), .B(n10408), .C(n10505), .Z(n10497) );
  HS65_LL_NAND4ABX3 U12668 ( .A(n10506), .B(n10364), .C(n10427), .D(n10497), 
        .Z(n10400) );
  HS65_LL_NOR4ABX2 U12669 ( .A(n10368), .B(n10367), .C(n10366), .D(n10365), 
        .Z(n10371) );
  HS65_LL_NOR4ABX2 U12670 ( .A(n10372), .B(n10371), .C(n10370), .D(n10369), 
        .Z(n10397) );
  HS65_LL_NOR2X2 U12671 ( .A(n10374), .B(n10373), .Z(n10471) );
  HS65_LL_NOR2X2 U12672 ( .A(n10410), .B(n10375), .Z(n15070) );
  HS65_LL_NOR4ABX2 U12673 ( .A(n10471), .B(n15070), .C(n10377), .D(n10376), 
        .Z(n10378) );
  HS65_LL_NAND3X2 U12674 ( .A(n15074), .B(n10379), .C(n10378), .Z(n10421) );
  HS65_LL_NAND4ABX3 U12675 ( .A(n10382), .B(n10421), .C(n10381), .D(n10380), 
        .Z(n10395) );
  HS65_LL_NAND2X2 U12676 ( .A(n10384), .B(n10383), .Z(n10426) );
  HS65_LL_NAND3AX3 U12677 ( .A(n10426), .B(n10386), .C(n10385), .Z(n15061) );
  HS65_LL_NOR2X2 U12678 ( .A(n10490), .B(n10407), .Z(n10388) );
  HS65_LL_NAND4ABX3 U12679 ( .A(n10469), .B(n10389), .C(n10388), .D(n10387), 
        .Z(n10393) );
  HS65_LL_NOR4ABX2 U12680 ( .A(n10471), .B(n10392), .C(n10391), .D(n10390), 
        .Z(n10518) );
  HS65_LL_NAND4ABX3 U12681 ( .A(n15061), .B(n10393), .C(n10497), .D(n10518), 
        .Z(n10394) );
  HS65_LL_AOI22X1 U12682 ( .A(n15088), .B(n10395), .C(n15084), .D(n10394), .Z(
        n10396) );
  HS65_LL_CBI4I1X3 U12683 ( .A(n10398), .B(n10397), .C(n10527), .D(n10396), 
        .Z(n10399) );
  HS65_LL_CBI4I6X2 U12684 ( .A(n10401), .B(n10400), .C(n15082), .D(n10399), 
        .Z(n10402) );
  HS65_LLS_XOR3X2 U12685 ( .A(n10402), .B(\u0/rcon [30]), .C(w0[30]), .Z(
        n15101) );
  HS65_LL_MUX21I1X3 U12686 ( .D0(n15101), .D1(key[126]), .S0(n11617), .Z(
        \u0/N72 ) );
  HS65_LL_MUX21I1X3 U12687 ( .D0(n10403), .D1(key[89]), .S0(n11617), .Z(
        \u0/N133 ) );
  HS65_LL_MUX21I1X3 U12688 ( .D0(n10404), .D1(key[45]), .S0(n11617), .Z(
        \u0/N187 ) );
  HS65_LL_MUX21I1X3 U12689 ( .D0(n14819), .D1(n14819), .S0(w0[2]), .Z(N479) );
  HS65_LL_NAND4ABX3 U12690 ( .A(n10407), .B(n10406), .C(n10504), .D(n10405), 
        .Z(n10440) );
  HS65_LL_NOR2X2 U12691 ( .A(n10521), .B(n10501), .Z(n10498) );
  HS65_LL_NAND4ABX3 U12692 ( .A(n10409), .B(n10408), .C(n10498), .D(n10512), 
        .Z(n10439) );
  HS65_LL_NOR2X2 U12693 ( .A(n10506), .B(n10410), .Z(n15060) );
  HS65_LL_NAND2X2 U12694 ( .A(n10412), .B(n10411), .Z(n15073) );
  HS65_LL_NAND4ABX3 U12695 ( .A(n15073), .B(n10415), .C(n10414), .D(n10413), 
        .Z(n10416) );
  HS65_LL_NOR4ABX2 U12696 ( .A(n15060), .B(n10418), .C(n10417), .D(n10416), 
        .Z(n10436) );
  HS65_LL_NOR2X2 U12697 ( .A(n10419), .B(n10502), .Z(n10451) );
  HS65_LL_AOI112X2 U12698 ( .A(n10423), .B(n10422), .C(n10421), .D(n10420), 
        .Z(n10424) );
  HS65_LL_NAND3X2 U12699 ( .A(n10425), .B(n10451), .C(n10424), .Z(n10433) );
  HS65_LL_NOR4ABX2 U12700 ( .A(n15070), .B(n10427), .C(n10521), .D(n10426), 
        .Z(n10429) );
  HS65_LL_NOR4ABX2 U12701 ( .A(n10504), .B(n10429), .C(n10456), .D(n10428), 
        .Z(n10430) );
  HS65_LL_AOI12X2 U12702 ( .A(n10431), .B(n10430), .C(n10527), .Z(n10432) );
  HS65_LL_CBI4I6X2 U12703 ( .A(n10434), .B(n10433), .C(n15084), .D(n10432), 
        .Z(n10435) );
  HS65_LL_CBI4I1X3 U12704 ( .A(n10437), .B(n10436), .C(n10535), .D(n10435), 
        .Z(n10438) );
  HS65_LL_CBI4I6X2 U12705 ( .A(n10440), .B(n10439), .C(n15088), .D(n10438), 
        .Z(n10441) );
  HS65_LLS_XOR3X2 U12706 ( .A(n10441), .B(\u0/rcon [24]), .C(w0[24]), .Z(
        n15103) );
  HS65_LL_MUX21I1X3 U12707 ( .D0(n15103), .D1(key[120]), .S0(n11617), .Z(
        \u0/N66 ) );
  HS65_LL_NAND4ABX3 U12708 ( .A(n10453), .B(n10443), .C(n10486), .D(n10442), 
        .Z(n10445) );
  HS65_LL_NAND4ABX3 U12709 ( .A(n15050), .B(n10445), .C(n10444), .D(n10518), 
        .Z(n10480) );
  HS65_LL_NAND2AX4 U12710 ( .A(n10492), .B(n10446), .Z(n15049) );
  HS65_LL_NAND4ABX3 U12711 ( .A(n10449), .B(n15049), .C(n10448), .D(n10447), 
        .Z(n10452) );
  HS65_LL_NAND4ABX3 U12712 ( .A(n10453), .B(n10452), .C(n10451), .D(n10450), 
        .Z(n10515) );
  HS65_LL_NOR4ABX2 U12713 ( .A(n10455), .B(n10454), .C(n15068), .D(n10515), 
        .Z(n10457) );
  HS65_LL_NOR4ABX2 U12714 ( .A(n10458), .B(n10457), .C(n10506), .D(n10456), 
        .Z(n10477) );
  HS65_LL_NOR4ABX2 U12715 ( .A(n10508), .B(n15075), .C(n10460), .D(n10459), 
        .Z(n10461) );
  HS65_LL_NAND4ABX3 U12716 ( .A(n10464), .B(n10463), .C(n10462), .D(n10461), 
        .Z(n10466) );
  HS65_LL_NAND4ABX3 U12717 ( .A(n10467), .B(n10466), .C(n10465), .D(n10537), 
        .Z(n10475) );
  HS65_LL_NOR2X2 U12718 ( .A(n10492), .B(n10468), .Z(n15064) );
  HS65_LL_NOR4ABX2 U12719 ( .A(n10471), .B(n10470), .C(n10496), .D(n10469), 
        .Z(n10472) );
  HS65_LL_NAND4ABX3 U12720 ( .A(n10490), .B(n10473), .C(n15064), .D(n10472), 
        .Z(n10474) );
  HS65_LL_AOI22X1 U12721 ( .A(n15082), .B(n10475), .C(n15088), .D(n10474), .Z(
        n10476) );
  HS65_LL_CBI4I1X3 U12722 ( .A(n10478), .B(n10477), .C(n10527), .D(n10476), 
        .Z(n10479) );
  HS65_LL_CBI4I6X2 U12723 ( .A(n10481), .B(n10480), .C(n15084), .D(n10479), 
        .Z(n10482) );
  HS65_LLS_XOR3X2 U12724 ( .A(n10482), .B(\u0/rcon [27]), .C(w0[27]), .Z(
        n15105) );
  HS65_LL_MUX21I1X3 U12725 ( .D0(n15105), .D1(key[123]), .S0(n15110), .Z(
        \u0/N69 ) );
  HS65_LL_MUX21I1X3 U12726 ( .D0(n10483), .D1(key[93]), .S0(n11617), .Z(
        \u0/N137 ) );
  HS65_LL_NOR4ABX2 U12727 ( .A(n10487), .B(n10486), .C(n10485), .D(n10484), 
        .Z(n10488) );
  HS65_LL_NAND3X2 U12728 ( .A(n10530), .B(n10488), .C(n10508), .Z(n15081) );
  HS65_LL_NAND2AX4 U12729 ( .A(n10490), .B(n10489), .Z(n10491) );
  HS65_LL_NOR3X1 U12730 ( .A(n10493), .B(n10492), .C(n10491), .Z(n10503) );
  HS65_LL_NAND4ABX3 U12731 ( .A(n10496), .B(n10495), .C(n10503), .D(n10494), 
        .Z(n10499) );
  HS65_LL_NAND4ABX3 U12732 ( .A(n10500), .B(n10499), .C(n10498), .D(n10497), 
        .Z(n10539) );
  HS65_LL_NOR4ABX2 U12733 ( .A(n10504), .B(n10503), .C(n10502), .D(n10501), 
        .Z(n10507) );
  HS65_LL_NOR4ABX2 U12734 ( .A(n10507), .B(n10528), .C(n10506), .D(n10505), 
        .Z(n10536) );
  HS65_LL_NAND4ABX3 U12735 ( .A(n10511), .B(n10510), .C(n10509), .D(n10508), 
        .Z(n10514) );
  HS65_LL_NAND4ABX3 U12736 ( .A(n10515), .B(n10514), .C(n10513), .D(n10512), 
        .Z(n10532) );
  HS65_LL_NAND3X2 U12737 ( .A(n10518), .B(n10517), .C(n10516), .Z(n10519) );
  HS65_LL_NOR3X1 U12738 ( .A(n10521), .B(n10520), .C(n10519), .Z(n15054) );
  HS65_LL_OAI21X2 U12739 ( .A(n10524), .B(n10523), .C(n10522), .Z(n10525) );
  HS65_LL_NOR4ABX2 U12740 ( .A(n15054), .B(n10526), .C(n15076), .D(n10525), 
        .Z(n10529) );
  HS65_LL_AOI13X2 U12741 ( .A(n10530), .B(n10529), .C(n10528), .D(n10527), .Z(
        n10531) );
  HS65_LL_CBI4I6X2 U12742 ( .A(n10533), .B(n10532), .C(n15088), .D(n10531), 
        .Z(n10534) );
  HS65_LL_CBI4I1X3 U12743 ( .A(n10537), .B(n10536), .C(n10535), .D(n10534), 
        .Z(n10538) );
  HS65_LL_CBI4I6X2 U12744 ( .A(n15081), .B(n10539), .C(n15084), .D(n10538), 
        .Z(n10540) );
  HS65_LLS_XOR3X2 U12745 ( .A(n10540), .B(\u0/rcon [26]), .C(w0[26]), .Z(
        n15107) );
  HS65_LL_MUX21I1X3 U12746 ( .D0(n15107), .D1(key[122]), .S0(n11617), .Z(
        \u0/N68 ) );
  HS65_LL_IVX2 U12747 ( .A(n15334), .Z(n15335) );
  HS65_LLS_XOR3X2 U12748 ( .A(n15510), .B(w2[26]), .C(n15192), .Z(n10541) );
  HS65_LL_MUXI21X2 U12749 ( .D0(n15334), .D1(n15335), .S0(n10541), .Z(n10545)
         );
  HS65_LL_BFX4 U12750 ( .A(n14808), .Z(n14832) );
  HS65_LL_OAI21X2 U12751 ( .A(n15630), .B(n10545), .C(n14832), .Z(n10544) );
  HS65_LL_AOI12X2 U12752 ( .A(w2[26]), .B(text_in_r[58]), .C(n14808), .Z(
        n10542) );
  HS65_LL_OAI21X2 U12753 ( .A(w2[26]), .B(text_in_r[58]), .C(n10542), .Z(
        n10543) );
  HS65_LL_CBI4I1X3 U12754 ( .A(n10545), .B(n15630), .C(n10544), .D(n10543), 
        .Z(N148) );
  HS65_LL_MUX21I1X3 U12755 ( .D0(n10546), .D1(key[57]), .S0(n11617), .Z(
        \u0/N199 ) );
  HS65_LL_NOR2X2 U12756 ( .A(n10552), .B(n14430), .Z(n10761) );
  HS65_LL_NOR2X2 U12757 ( .A(n10761), .B(n11577), .Z(n10571) );
  HS65_LL_NOR2X2 U12758 ( .A(n10547), .B(n11001), .Z(n11083) );
  HS65_LL_NOR2X2 U12759 ( .A(n10569), .B(n10567), .Z(n10793) );
  HS65_LL_NOR4ABX2 U12760 ( .A(n11083), .B(n10580), .C(n10793), .D(n11790), 
        .Z(n10548) );
  HS65_LL_NOR4ABX2 U12761 ( .A(n10571), .B(n10548), .C(n10589), .D(n10574), 
        .Z(n14444) );
  HS65_LL_NAND2X2 U12762 ( .A(n10553), .B(n10549), .Z(n14419) );
  HS65_LL_NAND3AX3 U12763 ( .A(n10562), .B(n10550), .C(n14419), .Z(n11580) );
  HS65_LL_NOR2X2 U12764 ( .A(n11573), .B(n10551), .Z(n11803) );
  HS65_LL_IVX2 U12765 ( .A(n10552), .Z(n10554) );
  HS65_LL_NAND2X2 U12766 ( .A(n10554), .B(n10553), .Z(n11789) );
  HS65_LL_NAND2X2 U12767 ( .A(n10555), .B(n14407), .Z(n10592) );
  HS65_LL_NOR4ABX2 U12768 ( .A(n11789), .B(n11574), .C(n10556), .D(n10592), 
        .Z(n10557) );
  HS65_LL_NAND3X2 U12769 ( .A(n10557), .B(n10599), .C(n10763), .Z(n11608) );
  HS65_LL_NOR2AX3 U12770 ( .A(n10558), .B(n11608), .Z(n11784) );
  HS65_LL_NAND4ABX3 U12771 ( .A(n11606), .B(n10559), .C(n11803), .D(n11784), 
        .Z(n10560) );
  HS65_LL_NOR4ABX2 U12772 ( .A(n14444), .B(n14432), .C(n11580), .D(n10560), 
        .Z(n10605) );
  HS65_LL_NAND2X2 U12773 ( .A(n10561), .B(n14407), .Z(n10776) );
  HS65_LL_NAND2AX4 U12774 ( .A(n14437), .B(n10599), .Z(n14425) );
  HS65_LL_NOR2X2 U12775 ( .A(n10563), .B(n10562), .Z(n10983) );
  HS65_LL_NOR2X2 U12776 ( .A(n10581), .B(n10979), .Z(n11002) );
  HS65_LL_NOR2AX3 U12777 ( .A(n10564), .B(sa01[0]), .Z(n10764) );
  HS65_LL_NOR2X2 U12778 ( .A(n10999), .B(n10764), .Z(n11600) );
  HS65_LL_NAND4ABX3 U12779 ( .A(n11606), .B(n10565), .C(n11002), .D(n11600), 
        .Z(n11787) );
  HS65_LL_IVX2 U12780 ( .A(n10566), .Z(n10568) );
  HS65_LL_NOR2X2 U12781 ( .A(n10762), .B(n10567), .Z(n11774) );
  HS65_LL_NOR2X2 U12782 ( .A(n11774), .B(n10982), .Z(n11799) );
  HS65_LL_OAI21X2 U12783 ( .A(n10569), .B(n10568), .C(n11799), .Z(n10570) );
  HS65_LL_NOR3X1 U12784 ( .A(n11793), .B(n11787), .C(n10570), .Z(n11082) );
  HS65_LL_NAND4ABX3 U12785 ( .A(n10776), .B(n14425), .C(n10983), .D(n11082), 
        .Z(n10588) );
  HS65_LL_NOR4ABX2 U12786 ( .A(n10571), .B(n10785), .C(n11074), .D(n11582), 
        .Z(n11785) );
  HS65_LL_NAND4ABX3 U12787 ( .A(n10778), .B(n11790), .C(n11785), .D(n11803), 
        .Z(n10587) );
  HS65_LL_NOR2X2 U12788 ( .A(n10573), .B(n10572), .Z(n10978) );
  HS65_LL_NOR2X2 U12789 ( .A(n10978), .B(n10574), .Z(n10977) );
  HS65_LL_IVX2 U12790 ( .A(n10987), .Z(n11090) );
  HS65_LL_AOI12X2 U12791 ( .A(n11090), .B(n10575), .C(n10982), .Z(n10576) );
  HS65_LL_NAND3X2 U12792 ( .A(n10977), .B(n10576), .C(n10763), .Z(n14414) );
  HS65_LL_NAND4ABX3 U12793 ( .A(n10578), .B(n11783), .C(n10787), .D(n10577), 
        .Z(n10579) );
  HS65_LL_NOR3AX2 U12794 ( .A(n10580), .B(n14414), .C(n10579), .Z(n11087) );
  HS65_LL_NOR2X2 U12795 ( .A(n10581), .B(n10778), .Z(n10582) );
  HS65_LL_NOR4ABX2 U12796 ( .A(n10582), .B(n14407), .C(n14438), .D(n10590), 
        .Z(n14417) );
  HS65_LL_NAND3X2 U12797 ( .A(sa01[7]), .B(sa01[6]), .C(n11091), .Z(n10773) );
  HS65_LL_NOR2X2 U12798 ( .A(n11606), .B(n10985), .Z(n10780) );
  HS65_LL_IVX2 U12799 ( .A(n10583), .Z(n10790) );
  HS65_LL_NAND2X2 U12800 ( .A(n10780), .B(n10790), .Z(n10996) );
  HS65_LL_NOR4ABX2 U12801 ( .A(n10773), .B(n10584), .C(n14424), .D(n10996), 
        .Z(n10585) );
  HS65_LL_AOI13X2 U12802 ( .A(n11087), .B(n14417), .C(n10585), .D(n11611), .Z(
        n10586) );
  HS65_LL_CBI4I6X2 U12803 ( .A(n10588), .B(n10587), .C(n14449), .D(n10586), 
        .Z(n10604) );
  HS65_LL_NOR3X1 U12804 ( .A(n10589), .B(n10979), .C(n11000), .Z(n11100) );
  HS65_LL_NAND4ABX3 U12805 ( .A(n11774), .B(n10590), .C(n11100), .D(n10787), 
        .Z(n10602) );
  HS65_LL_NAND4ABX3 U12806 ( .A(n11798), .B(n10592), .C(n10591), .D(n11792), 
        .Z(n10600) );
  HS65_LL_NOR2X2 U12807 ( .A(n10593), .B(n11573), .Z(n11781) );
  HS65_LL_NAND4ABX3 U12808 ( .A(n10596), .B(n10595), .C(n10594), .D(n14423), 
        .Z(n10597) );
  HS65_LL_NOR4ABX2 U12809 ( .A(n11781), .B(n10598), .C(n11606), .D(n10597), 
        .Z(n11017) );
  HS65_LL_NAND4ABX3 U12810 ( .A(n11577), .B(n10600), .C(n11017), .D(n10599), 
        .Z(n10601) );
  HS65_LL_OAI13X1 U12811 ( .A(n10602), .B(n10783), .C(n10601), .D(n14453), .Z(
        n10603) );
  HS65_LL_OAI112X1 U12812 ( .A(n10605), .B(n11587), .C(n10604), .D(n10603), 
        .Z(n15127) );
  HS65_LL_NOR3X1 U12813 ( .A(n10607), .B(n10711), .C(n10606), .Z(n10812) );
  HS65_LL_NOR4ABX2 U12814 ( .A(n10812), .B(n10626), .C(n10609), .D(n10608), 
        .Z(n10611) );
  HS65_LL_NOR3AX2 U12815 ( .A(n11056), .B(n13369), .C(n13378), .Z(n10610) );
  HS65_LL_NAND3X2 U12816 ( .A(n10820), .B(n10611), .C(n10610), .Z(n10652) );
  HS65_LL_NOR2X2 U12817 ( .A(n13366), .B(n11050), .Z(n10965) );
  HS65_LL_IVX2 U12818 ( .A(n10734), .Z(n10645) );
  HS65_LL_NAND2X2 U12819 ( .A(n10738), .B(n10645), .Z(n10967) );
  HS65_LL_OAI21X2 U12820 ( .A(n10957), .B(n10612), .C(n10956), .Z(n10949) );
  HS65_LL_NAND3AX3 U12821 ( .A(n10967), .B(n10944), .C(n10949), .Z(n13403) );
  HS65_LL_NOR4ABX2 U12822 ( .A(n10614), .B(n10613), .C(n10825), .D(n13403), 
        .Z(n10615) );
  HS65_LL_NAND4ABX3 U12823 ( .A(n10951), .B(n10616), .C(n10965), .D(n10615), 
        .Z(n11059) );
  HS65_LL_NOR4ABX2 U12824 ( .A(n10618), .B(n10617), .C(n10638), .D(n10715), 
        .Z(n13390) );
  HS65_LL_NAND4ABX3 U12825 ( .A(n10736), .B(n10619), .C(n11022), .D(n13390), 
        .Z(n10622) );
  HS65_LL_AOI12X2 U12826 ( .A(n10745), .B(sa12[6]), .C(n10620), .Z(n10718) );
  HS65_LL_NAND4ABX3 U12827 ( .A(n11059), .B(n10622), .C(n10718), .D(n10621), 
        .Z(n10651) );
  HS65_LL_IVX2 U12828 ( .A(n10756), .Z(n13393) );
  HS65_LL_NAND3X2 U12829 ( .A(sa12[1]), .B(n10741), .C(n10623), .Z(n10625) );
  HS65_LL_NOR4ABX2 U12830 ( .A(n10626), .B(n10625), .C(n13400), .D(n10624), 
        .Z(n10627) );
  HS65_LL_OAI112X1 U12831 ( .A(n10630), .B(n10629), .C(n10628), .D(n10627), 
        .Z(n10940) );
  HS65_LL_AND2X4 U12832 ( .A(n11057), .B(n10645), .Z(n10632) );
  HS65_LL_NOR4ABX2 U12833 ( .A(n10632), .B(n11030), .C(n10833), .D(n10631), 
        .Z(n10633) );
  HS65_LL_NAND4ABX3 U12834 ( .A(n10638), .B(n10940), .C(n10633), .D(n10735), 
        .Z(n10636) );
  HS65_LL_NOR3X1 U12835 ( .A(n10829), .B(n11051), .C(n10634), .Z(n10635) );
  HS65_LL_NAND4ABX3 U12836 ( .A(n10722), .B(n10636), .C(n10713), .D(n10635), 
        .Z(n10650) );
  HS65_LL_NAND4ABX3 U12837 ( .A(n10934), .B(n10638), .C(n10637), .D(n13367), 
        .Z(n10648) );
  HS65_LL_NAND4ABX3 U12838 ( .A(n10962), .B(n10639), .C(n10812), .D(n10963), 
        .Z(n10647) );
  HS65_LL_NOR4ABX2 U12839 ( .A(n10640), .B(n10948), .C(n11043), .D(n11050), 
        .Z(n10946) );
  HS65_LL_NOR2X2 U12840 ( .A(sa12[6]), .B(sa12[7]), .Z(n10642) );
  HS65_LL_NAND2X2 U12841 ( .A(n10642), .B(n10641), .Z(n10747) );
  HS65_LL_NOR4ABX2 U12842 ( .A(n10644), .B(n10732), .C(n10643), .D(n10950), 
        .Z(n10821) );
  HS65_LL_NAND3X2 U12843 ( .A(n10821), .B(n10645), .C(n10806), .Z(n10646) );
  HS65_LL_NOR3AX2 U12844 ( .A(n10747), .B(n11051), .C(n10646), .Z(n11039) );
  HS65_LL_NAND4ABX3 U12845 ( .A(n10648), .B(n10647), .C(n10946), .D(n11039), 
        .Z(n10649) );
  HS65_LL_MX41X4 U12846 ( .D0(n10652), .S0(n11068), .D1(n10651), .S1(n13393), 
        .D2(n10650), .S2(n13401), .D3(n10649), .S3(n13410), .Z(n15267) );
  HS65_LL_IVX2 U12847 ( .A(w1[30]), .Z(n15126) );
  HS65_LL_MUXI21X2 U12848 ( .D0(n15126), .D1(w1[30]), .S0(n15445), .Z(n10653)
         );
  HS65_LLS_XOR3X2 U12849 ( .A(n15127), .B(n15267), .C(n10653), .Z(n10710) );
  HS65_LL_NOR2X2 U12850 ( .A(n10859), .B(n14319), .Z(n11838) );
  HS65_LL_NOR2X2 U12851 ( .A(n11866), .B(n12213), .Z(n10668) );
  HS65_LL_NAND2X2 U12852 ( .A(n10660), .B(n10654), .Z(n13417) );
  HS65_LL_CBI4I1X3 U12853 ( .A(n10656), .B(n14309), .C(n10655), .D(n14296), 
        .Z(n10657) );
  HS65_LL_NOR4ABX2 U12854 ( .A(n10668), .B(n13417), .C(n11817), .D(n10657), 
        .Z(n14326) );
  HS65_LL_NAND2X2 U12855 ( .A(n10658), .B(n12202), .Z(n11828) );
  HS65_LL_NAND2X2 U12856 ( .A(n11828), .B(n11844), .Z(n10673) );
  HS65_LL_NAND2X2 U12857 ( .A(sa23[7]), .B(n10667), .Z(n10677) );
  HS65_LL_NAND2X2 U12858 ( .A(n11867), .B(n10677), .Z(n11883) );
  HS65_LL_NOR3X1 U12859 ( .A(n10687), .B(n10673), .C(n11883), .Z(n10876) );
  HS65_LL_NAND2X2 U12860 ( .A(n12201), .B(n10659), .Z(n14314) );
  HS65_LL_NAND2X2 U12861 ( .A(n14314), .B(n11841), .Z(n11832) );
  HS65_LL_NOR4ABX2 U12862 ( .A(n14326), .B(n10876), .C(n12220), .D(n11832), 
        .Z(n10663) );
  HS65_LL_IVX2 U12863 ( .A(n14299), .Z(n13431) );
  HS65_LL_NAND2X2 U12864 ( .A(n10660), .B(n12202), .Z(n11840) );
  HS65_LL_NAND3X2 U12865 ( .A(n13431), .B(n11840), .C(n12196), .Z(n11826) );
  HS65_LL_NAND2X2 U12866 ( .A(n10661), .B(n10671), .Z(n13414) );
  HS65_LL_NAND3AX3 U12867 ( .A(n13414), .B(n10697), .C(n11825), .Z(n11879) );
  HS65_LL_NOR2X2 U12868 ( .A(n13452), .B(n14328), .Z(n12210) );
  HS65_LL_OAI21X2 U12869 ( .A(n14317), .B(n10664), .C(n11872), .Z(n13445) );
  HS65_LL_NOR4ABX2 U12870 ( .A(n12210), .B(n11845), .C(n11827), .D(n13445), 
        .Z(n10662) );
  HS65_LL_NAND4ABX3 U12871 ( .A(n14291), .B(n11879), .C(n10662), .D(n10698), 
        .Z(n10858) );
  HS65_LL_NOR4ABX2 U12872 ( .A(n11838), .B(n10663), .C(n11826), .D(n10858), 
        .Z(n10706) );
  HS65_LL_NOR3X1 U12873 ( .A(n10666), .B(n10665), .C(n10664), .Z(n13437) );
  HS65_LL_NAND3AX3 U12874 ( .A(n13437), .B(n10698), .C(n11828), .Z(n12226) );
  HS65_LL_OR2X4 U12875 ( .A(n10667), .B(n13422), .Z(n10864) );
  HS65_LL_NOR4ABX2 U12876 ( .A(n11882), .B(n10668), .C(n12226), .D(n10864), 
        .Z(n10669) );
  HS65_LL_NAND3X2 U12877 ( .A(n10669), .B(n11860), .C(n11833), .Z(n11847) );
  HS65_LL_NAND2X2 U12878 ( .A(n10670), .B(n11816), .Z(n11878) );
  HS65_LL_NAND4ABX3 U12879 ( .A(n11878), .B(n10672), .C(n10671), .D(n14296), 
        .Z(n10686) );
  HS65_LL_NOR2X2 U12880 ( .A(n10674), .B(n10673), .Z(n11890) );
  HS65_LL_NOR3X1 U12881 ( .A(n10675), .B(n14291), .C(n13414), .Z(n10846) );
  HS65_LL_NOR2X2 U12882 ( .A(sa23[5]), .B(n10676), .Z(n14304) );
  HS65_LL_NOR2X2 U12883 ( .A(n11827), .B(n14304), .Z(n11834) );
  HS65_LL_NAND2AX4 U12884 ( .A(n13422), .B(n10697), .Z(n13421) );
  HS65_LL_NAND3X2 U12885 ( .A(n10678), .B(n11815), .C(n10677), .Z(n10679) );
  HS65_LL_NOR3X1 U12886 ( .A(n10680), .B(n13421), .C(n10679), .Z(n13453) );
  HS65_LL_NAND2X2 U12887 ( .A(n10681), .B(n10851), .Z(n14320) );
  HS65_LL_IVX2 U12888 ( .A(n14320), .Z(n10855) );
  HS65_LL_NOR2X2 U12889 ( .A(n10855), .B(n10682), .Z(n11842) );
  HS65_LL_NAND2X2 U12890 ( .A(n11842), .B(n11816), .Z(n12207) );
  HS65_LL_NAND4ABX3 U12891 ( .A(n13452), .B(n13438), .C(n14326), .D(n13423), 
        .Z(n10683) );
  HS65_LL_NOR4ABX2 U12892 ( .A(n11834), .B(n13453), .C(n12207), .D(n10683), 
        .Z(n10684) );
  HS65_LL_AOI13X2 U12893 ( .A(n11890), .B(n10846), .C(n10684), .D(n12229), .Z(
        n10685) );
  HS65_LL_CBI4I6X2 U12894 ( .A(n11847), .B(n10686), .C(n14337), .D(n10685), 
        .Z(n10705) );
  HS65_LL_IVX2 U12895 ( .A(n10687), .Z(n11874) );
  HS65_LL_NAND4ABX3 U12896 ( .A(n11817), .B(n12200), .C(n10688), .D(n11874), 
        .Z(n10703) );
  HS65_LL_NAND2X2 U12897 ( .A(n10689), .B(n13448), .Z(n11855) );
  HS65_LL_NOR2X2 U12898 ( .A(n11863), .B(n10690), .Z(n13416) );
  HS65_LL_NOR2X2 U12899 ( .A(n10691), .B(n13416), .Z(n10863) );
  HS65_LL_NOR4ABX2 U12900 ( .A(n10863), .B(n10693), .C(n10692), .D(n13438), 
        .Z(n10694) );
  HS65_LL_NAND4ABX3 U12901 ( .A(n11855), .B(n13456), .C(n11842), .D(n10694), 
        .Z(n12195) );
  HS65_LL_IVX2 U12902 ( .A(n11841), .Z(n10865) );
  HS65_LL_NOR2X2 U12903 ( .A(n10865), .B(n14319), .Z(n11873) );
  HS65_LL_AND2X4 U12904 ( .A(n10695), .B(n11873), .Z(n13418) );
  HS65_LL_NAND2X2 U12905 ( .A(n10696), .B(n10852), .Z(n12203) );
  HS65_LL_NAND2X2 U12906 ( .A(n10697), .B(n12203), .Z(n11848) );
  HS65_LL_NAND4ABX3 U12907 ( .A(n12220), .B(n11848), .C(n10698), .D(n14296), 
        .Z(n10699) );
  HS65_LL_AOI12X2 U12908 ( .A(n10700), .B(n12201), .C(n10699), .Z(n10848) );
  HS65_LL_NAND4ABX3 U12909 ( .A(n10859), .B(n10701), .C(n13418), .D(n10848), 
        .Z(n10702) );
  HS65_LL_OAI13X1 U12910 ( .A(n10703), .B(n12195), .C(n10702), .D(n14335), .Z(
        n10704) );
  HS65_LL_OAI112X1 U12911 ( .A(n10706), .B(n11880), .C(n10705), .D(n10704), 
        .Z(n14955) );
  HS65_LL_IVX2 U12912 ( .A(n14955), .Z(n15359) );
  HS65_LL_MUXI21X2 U12913 ( .D0(n14955), .D1(n15359), .S0(n15266), .Z(n14544)
         );
  HS65_LL_OAI21X2 U12914 ( .A(n14544), .B(n10710), .C(n14832), .Z(n10709) );
  HS65_LL_IVX2 U12915 ( .A(text_in_r[94]), .Z(n10707) );
  HS65_LL_IVX4 U12916 ( .A(n11557), .Z(n15545) );
  HS65_LL_OAI212X3 U12917 ( .A(w1[30]), .B(text_in_r[94]), .C(n15126), .D(
        n10707), .E(n15545), .Z(n10708) );
  HS65_LL_CBI4I1X3 U12918 ( .A(n10710), .B(n14544), .C(n10709), .D(n10708), 
        .Z(N216) );
  HS65_LL_IVX4 U12919 ( .A(n14808), .Z(n15688) );
  HS65_LL_OAI21X2 U12920 ( .A(w1[25]), .B(text_in_r[89]), .C(n15688), .Z(
        n11021) );
  HS65_LL_IVX2 U12921 ( .A(n11557), .Z(n14822) );
  HS65_LL_NOR4ABX2 U12922 ( .A(n10713), .B(n10712), .C(n10711), .D(n13377), 
        .Z(n10714) );
  HS65_LL_NAND4ABX3 U12923 ( .A(n10716), .B(n10715), .C(n11031), .D(n10714), 
        .Z(n10760) );
  HS65_LL_NAND2X2 U12924 ( .A(n10717), .B(n11052), .Z(n13376) );
  HS65_LL_OAI21X2 U12925 ( .A(n10720), .B(n10719), .C(n10718), .Z(n10721) );
  HS65_LL_NOR3X1 U12926 ( .A(n10722), .B(n13376), .C(n10721), .Z(n11040) );
  HS65_LL_NOR4ABX2 U12927 ( .A(n10821), .B(n10724), .C(n10934), .D(n10723), 
        .Z(n10727) );
  HS65_LL_NAND2X2 U12928 ( .A(n10726), .B(n10725), .Z(n13399) );
  HS65_LL_NOR4ABX2 U12929 ( .A(n11040), .B(n10727), .C(n13382), .D(n13399), 
        .Z(n10757) );
  HS65_LL_NAND2X2 U12930 ( .A(n10728), .B(n11041), .Z(n10832) );
  HS65_LL_NOR4ABX2 U12931 ( .A(n10731), .B(n10730), .C(n10729), .D(n10832), 
        .Z(n10733) );
  HS65_LL_NAND4ABX3 U12932 ( .A(n10734), .B(n13369), .C(n10733), .D(n10732), 
        .Z(n10753) );
  HS65_LL_NOR2X2 U12933 ( .A(n13366), .B(n13400), .Z(n10816) );
  HS65_LL_NAND4ABX3 U12934 ( .A(n10736), .B(n13377), .C(n10816), .D(n10735), 
        .Z(n10737) );
  HS65_LL_NOR3X1 U12935 ( .A(n10962), .B(n13365), .C(n10737), .Z(n10836) );
  HS65_LL_NAND2X2 U12936 ( .A(n10739), .B(n10738), .Z(n10935) );
  HS65_LL_AOI12X2 U12937 ( .A(n10741), .B(n10740), .C(n10951), .Z(n11027) );
  HS65_LL_NAND3AX3 U12938 ( .A(n10743), .B(n11027), .C(n10742), .Z(n10744) );
  HS65_LL_NOR3X1 U12939 ( .A(n10811), .B(n10935), .C(n10744), .Z(n10818) );
  HS65_LL_NOR2X2 U12940 ( .A(n11043), .B(n13383), .Z(n10933) );
  HS65_LL_IVX2 U12941 ( .A(n10745), .Z(n10748) );
  HS65_LL_CBI4I1X3 U12942 ( .A(n10748), .B(n10747), .C(sa12[1]), .D(n10746), 
        .Z(n10749) );
  HS65_LL_NOR4ABX2 U12943 ( .A(n11031), .B(n10933), .C(n10934), .D(n10749), 
        .Z(n10751) );
  HS65_LL_AOI13X2 U12944 ( .A(n10836), .B(n10818), .C(n10751), .D(n10750), .Z(
        n10752) );
  HS65_LL_CBI4I6X2 U12945 ( .A(n10754), .B(n10753), .C(n13401), .D(n10752), 
        .Z(n10755) );
  HS65_LL_OAI21X2 U12946 ( .A(n10757), .B(n10756), .C(n10755), .Z(n10758) );
  HS65_LL_CBI4I6X2 U12947 ( .A(n10760), .B(n10759), .C(n11068), .D(n10758), 
        .Z(n15264) );
  HS65_LL_IVX2 U12948 ( .A(n15264), .Z(n15263) );
  HS65_LL_NOR2X2 U12949 ( .A(n10761), .B(n11774), .Z(n11594) );
  HS65_LL_OAI112X1 U12950 ( .A(n10762), .B(n10987), .C(n11594), .D(n14432), 
        .Z(n10804) );
  HS65_LL_NOR2X2 U12951 ( .A(n11601), .B(n14430), .Z(n11070) );
  HS65_LL_IVX2 U12952 ( .A(n10763), .Z(n11794) );
  HS65_LL_NOR2X2 U12953 ( .A(n10764), .B(n11794), .Z(n11005) );
  HS65_LL_AOI12X2 U12954 ( .A(n11078), .B(n10766), .C(n10765), .Z(n10767) );
  HS65_LL_NOR4ABX2 U12955 ( .A(n14433), .B(n10767), .C(n10999), .D(n11580), 
        .Z(n11570) );
  HS65_LL_NAND4ABX3 U12956 ( .A(n11070), .B(n14442), .C(n11005), .D(n11570), 
        .Z(n10769) );
  HS65_LL_NAND4ABX3 U12957 ( .A(n11597), .B(n10769), .C(n10768), .D(n14407), 
        .Z(n10803) );
  HS65_LL_NAND2X2 U12958 ( .A(n10771), .B(n10770), .Z(n10772) );
  HS65_LL_NAND2X2 U12959 ( .A(n11789), .B(n11802), .Z(n14441) );
  HS65_LL_NOR4ABX2 U12960 ( .A(n10773), .B(n10772), .C(n10798), .D(n14441), 
        .Z(n10994) );
  HS65_LL_NAND4ABX3 U12961 ( .A(n11787), .B(n10774), .C(n10974), .D(n14412), 
        .Z(n10775) );
  HS65_LL_NOR4ABX2 U12962 ( .A(n10994), .B(n14443), .C(n10776), .D(n10775), 
        .Z(n10801) );
  HS65_LL_NOR2X2 U12963 ( .A(n10777), .B(n10793), .Z(n11565) );
  HS65_LL_IVX2 U12964 ( .A(n10978), .Z(n10789) );
  HS65_LL_NOR4ABX2 U12965 ( .A(n10992), .B(n10789), .C(n10778), .D(n11805), 
        .Z(n10779) );
  HS65_LL_NAND4ABX3 U12966 ( .A(n14442), .B(n11790), .C(n11565), .D(n10779), 
        .Z(n11592) );
  HS65_LL_NAND2X2 U12967 ( .A(n10986), .B(n14408), .Z(n10995) );
  HS65_LL_NAND3X2 U12968 ( .A(n10780), .B(n11789), .C(n14407), .Z(n11569) );
  HS65_LL_NAND4ABX3 U12969 ( .A(n10995), .B(n11569), .C(n11083), .D(n10781), 
        .Z(n10782) );
  HS65_LL_OAI13X1 U12970 ( .A(n11592), .B(n10783), .C(n10782), .D(n14447), .Z(
        n10800) );
  HS65_LL_NOR2X2 U12971 ( .A(n10784), .B(n14438), .Z(n10998) );
  HS65_LL_NAND2X2 U12972 ( .A(n10998), .B(n10785), .Z(n10975) );
  HS65_LL_NAND2X2 U12973 ( .A(n10786), .B(n11574), .Z(n14410) );
  HS65_LL_NOR4ABX2 U12974 ( .A(n10983), .B(n14423), .C(n14424), .D(n11577), 
        .Z(n10788) );
  HS65_LL_NAND4ABX3 U12975 ( .A(n11783), .B(n14410), .C(n10788), .D(n10787), 
        .Z(n11809) );
  HS65_LL_NOR4ABX2 U12976 ( .A(n10789), .B(n14419), .C(n11805), .D(n11000), 
        .Z(n10791) );
  HS65_LL_NAND3X2 U12977 ( .A(n10792), .B(n10791), .C(n10790), .Z(n11782) );
  HS65_LL_IVX2 U12978 ( .A(n10793), .Z(n11788) );
  HS65_LL_NOR2X2 U12979 ( .A(sa01[1]), .B(n10794), .Z(n10795) );
  HS65_LL_AOI12X2 U12980 ( .A(n10795), .B(n11091), .C(n11569), .Z(n10796) );
  HS65_LL_NAND4ABX3 U12981 ( .A(n11809), .B(n11782), .C(n11788), .D(n10796), 
        .Z(n10797) );
  HS65_LL_OAI13X1 U12982 ( .A(n10798), .B(n10975), .C(n10797), .D(n14449), .Z(
        n10799) );
  HS65_LL_OAI112X1 U12983 ( .A(n10801), .B(n11611), .C(n10800), .D(n10799), 
        .Z(n10802) );
  HS65_LL_CBI4I6X2 U12984 ( .A(n10804), .B(n10803), .C(n14453), .D(n10802), 
        .Z(n15124) );
  HS65_LL_MUXI21X2 U12985 ( .D0(n15264), .D1(n15263), .S0(n15124), .Z(n10805)
         );
  HS65_LL_NOR2X2 U12986 ( .A(n14822), .B(n10805), .Z(n14842) );
  HS65_LL_IVX4 U12987 ( .A(n14808), .Z(n15698) );
  HS65_LL_NOR2AX3 U12988 ( .A(n10805), .B(n15698), .Z(n14843) );
  HS65_LL_NAND4ABX3 U12989 ( .A(n10951), .B(n13386), .C(n10807), .D(n10806), 
        .Z(n10808) );
  HS65_LL_AOI12X2 U12990 ( .A(n10810), .B(n10809), .C(n10808), .Z(n10947) );
  HS65_LL_NAND4ABX3 U12991 ( .A(n10811), .B(n10936), .C(n10947), .D(n11052), 
        .Z(n10813) );
  HS65_LL_NAND4ABX3 U12992 ( .A(n10814), .B(n10813), .C(n10836), .D(n10812), 
        .Z(n10841) );
  HS65_LL_NAND3X2 U12993 ( .A(n10816), .B(n10822), .C(n10815), .Z(n10817) );
  HS65_LL_NOR4ABX2 U12994 ( .A(n10818), .B(n10946), .C(n10930), .D(n10817), 
        .Z(n10819) );
  HS65_LL_NAND3X2 U12995 ( .A(n10821), .B(n10820), .C(n10819), .Z(n10840) );
  HS65_LL_NAND2X2 U12996 ( .A(n10823), .B(n10822), .Z(n13395) );
  HS65_LL_NOR2X2 U12997 ( .A(sa12[3]), .B(n10824), .Z(n10937) );
  HS65_LL_NAND4ABX3 U12998 ( .A(n10937), .B(n13382), .C(n11040), .D(n13372), 
        .Z(n10828) );
  HS65_LL_NOR3X1 U12999 ( .A(n10955), .B(n10825), .C(n11051), .Z(n10827) );
  HS65_LL_NAND4ABX3 U13000 ( .A(n13395), .B(n10828), .C(n10827), .D(n10826), 
        .Z(n10839) );
  HS65_LL_NOR4ABX2 U13001 ( .A(n10949), .B(n10948), .C(n13388), .D(n10829), 
        .Z(n10830) );
  HS65_LL_NAND4ABX3 U13002 ( .A(n11044), .B(n10832), .C(n10831), .D(n10830), 
        .Z(n13412) );
  HS65_LL_NOR4ABX2 U13003 ( .A(n10834), .B(n11030), .C(n10833), .D(n10967), 
        .Z(n10835) );
  HS65_LL_NAND4ABX3 U13004 ( .A(n10837), .B(n13412), .C(n10836), .D(n10835), 
        .Z(n10838) );
  HS65_LL_MX41X4 U13005 ( .D0(n10841), .S0(n11068), .D1(n10840), .S1(n13393), 
        .D2(n10839), .S2(n13401), .D3(n10838), .S3(n13410), .Z(n15273) );
  HS65_LL_OAI21X2 U13006 ( .A(n10842), .B(n11864), .C(n11815), .Z(n10843) );
  HS65_LL_NOR3X1 U13007 ( .A(n14299), .B(n10844), .C(n10843), .Z(n11836) );
  HS65_LL_NOR3X1 U13008 ( .A(n13451), .B(n13422), .C(n11832), .Z(n10845) );
  HS65_LL_NAND3X2 U13009 ( .A(n10846), .B(n10845), .C(n12197), .Z(n11858) );
  HS65_LL_NAND3X2 U13010 ( .A(n11840), .B(n13417), .C(n11872), .Z(n10847) );
  HS65_LL_NOR4ABX2 U13011 ( .A(n10848), .B(n10869), .C(n11858), .D(n10847), 
        .Z(n10849) );
  HS65_LL_NAND3X2 U13012 ( .A(n11836), .B(n10850), .C(n10849), .Z(n10880) );
  HS65_LL_IVX2 U13013 ( .A(n11880), .Z(n14339) );
  HS65_LL_AOI12X2 U13014 ( .A(n10852), .B(n10851), .C(n13428), .Z(n12199) );
  HS65_LL_NAND2X2 U13015 ( .A(n10874), .B(n12202), .Z(n10853) );
  HS65_LL_NAND3X2 U13016 ( .A(n12199), .B(n10853), .C(n13417), .Z(n10854) );
  HS65_LL_NOR3X1 U13017 ( .A(n13446), .B(n11855), .C(n10854), .Z(n11814) );
  HS65_LL_NAND2X2 U13018 ( .A(n11814), .B(n13418), .Z(n11885) );
  HS65_LL_AOI12X2 U13019 ( .A(n10857), .B(n10856), .C(n10855), .Z(n11829) );
  HS65_LL_NOR2X2 U13020 ( .A(n14292), .B(n10858), .Z(n13442) );
  HS65_LL_NOR4ABX2 U13021 ( .A(n11829), .B(n13442), .C(n10868), .D(n10859), 
        .Z(n10860) );
  HS65_LL_NAND4ABX3 U13022 ( .A(n13429), .B(n11885), .C(n10861), .D(n10860), 
        .Z(n10879) );
  HS65_LL_NAND2X2 U13023 ( .A(n10862), .B(n12197), .Z(n11835) );
  HS65_LL_NAND2X2 U13024 ( .A(n10863), .B(n11875), .Z(n11824) );
  HS65_LL_NOR3X1 U13025 ( .A(n14292), .B(n11824), .C(n10864), .Z(n10866) );
  HS65_LL_NAND4ABX3 U13026 ( .A(n11818), .B(n13432), .C(n11872), .D(n11815), 
        .Z(n11857) );
  HS65_LL_NOR4ABX2 U13027 ( .A(n10866), .B(n11828), .C(n10865), .D(n11857), 
        .Z(n10867) );
  HS65_LL_NAND4ABX3 U13028 ( .A(n11835), .B(n14313), .C(n11887), .D(n10867), 
        .Z(n10878) );
  HS65_LL_NOR2X2 U13029 ( .A(n11817), .B(n13433), .Z(n14323) );
  HS65_LL_NOR2X2 U13030 ( .A(n10868), .B(n13416), .Z(n11876) );
  HS65_LL_NAND3X2 U13031 ( .A(n12199), .B(n11876), .C(n10869), .Z(n10870) );
  HS65_LL_NOR3AX2 U13032 ( .A(n14323), .B(n10871), .C(n10870), .Z(n13450) );
  HS65_LL_NAND3X2 U13033 ( .A(n13436), .B(n11845), .C(n13423), .Z(n10872) );
  HS65_LL_AOI112X2 U13034 ( .A(n10874), .B(n10873), .C(n11858), .D(n10872), 
        .Z(n10875) );
  HS65_LL_NAND3X2 U13035 ( .A(n10876), .B(n13450), .C(n10875), .Z(n10877) );
  HS65_LL_MX41X4 U13036 ( .D0(n10880), .S0(n14339), .D1(n10879), .S1(n14337), 
        .D2(n10878), .S2(n14335), .D3(n10877), .S3(n14333), .Z(n15369) );
  HS65_LLS_XOR2X3 U13037 ( .A(n15273), .B(n15369), .Z(n14968) );
  HS65_LL_NOR4ABX2 U13038 ( .A(n12184), .B(n12835), .C(n12846), .D(n10881), 
        .Z(n10888) );
  HS65_LL_NAND3X2 U13039 ( .A(n10923), .B(n12173), .C(n10882), .Z(n10884) );
  HS65_LL_NAND4ABX3 U13040 ( .A(n10885), .B(n10884), .C(n12836), .D(n10883), 
        .Z(n11122) );
  HS65_LL_NOR3X1 U13041 ( .A(n12823), .B(n10886), .C(n11122), .Z(n10887) );
  HS65_LL_NAND3X2 U13042 ( .A(n11112), .B(n10888), .C(n10887), .Z(n10929) );
  HS65_LL_IVX2 U13043 ( .A(n11125), .Z(n10905) );
  HS65_LL_NAND2X2 U13044 ( .A(n11118), .B(n10905), .Z(n10891) );
  HS65_LL_NAND4ABX3 U13045 ( .A(n10891), .B(n10890), .C(n12169), .D(n10889), 
        .Z(n10892) );
  HS65_LL_NOR2X2 U13046 ( .A(n14657), .B(n11130), .Z(n14666) );
  HS65_LL_NAND4ABX3 U13047 ( .A(n10893), .B(n10892), .C(n14666), .D(n12829), 
        .Z(n14693) );
  HS65_LL_NOR4ABX2 U13048 ( .A(n10895), .B(n10894), .C(n12846), .D(n12176), 
        .Z(n10896) );
  HS65_LL_NAND3X2 U13049 ( .A(n10898), .B(n10897), .C(n10896), .Z(n11116) );
  HS65_LL_NOR4ABX2 U13050 ( .A(n10902), .B(n10901), .C(n10900), .D(n10899), 
        .Z(n10903) );
  HS65_LL_NAND4ABX3 U13051 ( .A(n14693), .B(n11116), .C(n10904), .D(n10903), 
        .Z(n10928) );
  HS65_LL_NAND2X2 U13052 ( .A(n10906), .B(n10905), .Z(n10914) );
  HS65_LL_NOR2X2 U13053 ( .A(sa30[1]), .B(n10907), .Z(n11115) );
  HS65_LL_OAI13X1 U13054 ( .A(sa30[6]), .B(n11115), .C(n10908), .D(n11113), 
        .Z(n10913) );
  HS65_LL_NOR4ABX2 U13055 ( .A(n11119), .B(n12174), .C(n14657), .D(n11131), 
        .Z(n10910) );
  HS65_LL_NAND3X2 U13056 ( .A(n10910), .B(n10909), .C(n12162), .Z(n12820) );
  HS65_LL_IVX2 U13057 ( .A(n12820), .Z(n11110) );
  HS65_LL_NOR4ABX2 U13058 ( .A(n14663), .B(n12850), .C(n10911), .D(n14648), 
        .Z(n10912) );
  HS65_LL_NAND4ABX3 U13059 ( .A(n10914), .B(n10913), .C(n11110), .D(n10912), 
        .Z(n10927) );
  HS65_LL_NAND3X2 U13060 ( .A(n10917), .B(n10916), .C(n10915), .Z(n10918) );
  HS65_LL_NOR3X1 U13061 ( .A(n10920), .B(n10919), .C(n10918), .Z(n12822) );
  HS65_LL_NOR4ABX2 U13062 ( .A(n10923), .B(n12162), .C(n10922), .D(n10921), 
        .Z(n10924) );
  HS65_LL_NAND4ABX3 U13063 ( .A(n11116), .B(n10925), .C(n12822), .D(n10924), 
        .Z(n10926) );
  HS65_LL_MX41X4 U13064 ( .D0(n10929), .S0(n12192), .D1(n10928), .S1(n14691), 
        .D2(n10927), .S2(n14683), .D3(n10926), .S3(n14685), .Z(n15451) );
  HS65_LL_NOR3X1 U13065 ( .A(n10931), .B(n10930), .C(n13375), .Z(n10932) );
  HS65_LL_NAND4ABX3 U13066 ( .A(n10934), .B(n13386), .C(n10933), .D(n10932), 
        .Z(n10939) );
  HS65_LL_NOR3X1 U13067 ( .A(n10937), .B(n10936), .C(n10935), .Z(n10938) );
  HS65_LL_NAND4ABX3 U13068 ( .A(n10940), .B(n10939), .C(n11040), .D(n10938), 
        .Z(n10971) );
  HS65_LL_NAND3X2 U13069 ( .A(n11056), .B(n10941), .C(n11045), .Z(n10942) );
  HS65_LL_NOR4ABX2 U13070 ( .A(n10944), .B(n10943), .C(n10950), .D(n10942), 
        .Z(n10945) );
  HS65_LL_NAND3X2 U13071 ( .A(n10947), .B(n10946), .C(n10945), .Z(n10970) );
  HS65_LL_NAND4ABX3 U13072 ( .A(n10951), .B(n10950), .C(n10949), .D(n10948), 
        .Z(n10953) );
  HS65_LL_NOR4ABX2 U13073 ( .A(n11056), .B(n11062), .C(n11064), .D(n13377), 
        .Z(n10952) );
  HS65_LL_NAND4ABX3 U13074 ( .A(n10954), .B(n10953), .C(n11040), .D(n10952), 
        .Z(n10969) );
  HS65_LL_AOI12X2 U13075 ( .A(n10957), .B(n10956), .C(n10955), .Z(n11026) );
  HS65_LL_NAND2X2 U13076 ( .A(sa12[7]), .B(n13392), .Z(n10959) );
  HS65_LL_AOI12X2 U13077 ( .A(n10960), .B(n10959), .C(n10958), .Z(n10961) );
  HS65_LL_NOR4ABX2 U13078 ( .A(n11026), .B(n10963), .C(n10962), .D(n10961), 
        .Z(n10964) );
  HS65_LL_NAND4ABX3 U13079 ( .A(n10967), .B(n10966), .C(n10965), .D(n10964), 
        .Z(n10968) );
  HS65_LL_MX41X4 U13080 ( .D0(n10971), .S0(n11068), .D1(n10970), .S1(n13393), 
        .D2(n10969), .S2(n13401), .D3(n10968), .S3(n13410), .Z(n15275) );
  HS65_LLS_XOR3X2 U13081 ( .A(w1[25]), .B(n15451), .C(n15275), .Z(n11018) );
  HS65_LL_NAND2X2 U13082 ( .A(n10994), .B(n10980), .Z(n11086) );
  HS65_LL_AOI12X2 U13083 ( .A(n10973), .B(n10972), .C(n11086), .Z(n11778) );
  HS65_LL_NAND4ABX3 U13084 ( .A(n10975), .B(n11804), .C(n11778), .D(n10974), 
        .Z(n10976) );
  HS65_LL_NOR4ABX2 U13085 ( .A(n10977), .B(n11780), .C(n14442), .D(n10976), 
        .Z(n11016) );
  HS65_LL_NOR2X2 U13086 ( .A(n10979), .B(n10978), .Z(n11593) );
  HS65_LL_AND2X4 U13087 ( .A(n11004), .B(n10980), .Z(n11095) );
  HS65_LL_NOR4ABX2 U13088 ( .A(n10983), .B(n11095), .C(n10982), .D(n10981), 
        .Z(n10984) );
  HS65_LL_NAND4ABX3 U13089 ( .A(n11783), .B(n10985), .C(n11593), .D(n10984), 
        .Z(n11013) );
  HS65_LL_OAI112X1 U13090 ( .A(n10988), .B(n10987), .C(n11586), .D(n10986), 
        .Z(n10989) );
  HS65_LL_NOR3X1 U13091 ( .A(n11000), .B(n11793), .C(n10989), .Z(n11807) );
  HS65_LL_NOR4ABX2 U13092 ( .A(n10992), .B(n11092), .C(n10991), .D(n10990), 
        .Z(n10993) );
  HS65_LL_NAND2X2 U13093 ( .A(n11002), .B(n14423), .Z(n11585) );
  HS65_LL_NOR4ABX2 U13094 ( .A(n11807), .B(n10993), .C(n11580), .D(n11585), 
        .Z(n11011) );
  HS65_LL_IVX2 U13095 ( .A(n10994), .Z(n11009) );
  HS65_LL_NOR3X1 U13096 ( .A(n10996), .B(n10995), .C(n14446), .Z(n10997) );
  HS65_LL_NAND4ABX3 U13097 ( .A(n11774), .B(n10999), .C(n10998), .D(n10997), 
        .Z(n11572) );
  HS65_LL_NOR2X2 U13098 ( .A(n11001), .B(n11000), .Z(n11604) );
  HS65_LL_NAND4ABX3 U13099 ( .A(n11580), .B(n11003), .C(n11002), .D(n11604), 
        .Z(n11006) );
  HS65_LL_NAND4ABX3 U13100 ( .A(n11007), .B(n11006), .C(n11005), .D(n11004), 
        .Z(n11008) );
  HS65_LL_OAI13X1 U13101 ( .A(n11009), .B(n11572), .C(n11008), .D(n14453), .Z(
        n11010) );
  HS65_LL_CBI4I1X3 U13102 ( .A(n11785), .B(n11011), .C(n11611), .D(n11010), 
        .Z(n11012) );
  HS65_LL_CBI4I6X2 U13103 ( .A(n11014), .B(n11013), .C(n14449), .D(n11012), 
        .Z(n11015) );
  HS65_LL_CBI4I1X3 U13104 ( .A(n11017), .B(n11016), .C(n11587), .D(n11015), 
        .Z(n15137) );
  HS65_LLS_XOR3X2 U13105 ( .A(n14968), .B(n11018), .C(n15137), .Z(n11019) );
  HS65_LL_MUXI21X2 U13106 ( .D0(n14842), .D1(n14843), .S0(n11019), .Z(n11020)
         );
  HS65_LL_CBI4I1X3 U13107 ( .A(text_in_r[89]), .B(w1[25]), .C(n11021), .D(
        n11020), .Z(N211) );
  HS65_LL_OAI112X1 U13108 ( .A(n11025), .B(n11024), .C(n11023), .D(n11022), 
        .Z(n11029) );
  HS65_LL_NOR4ABX2 U13109 ( .A(n11027), .B(n11026), .C(n11048), .D(n13387), 
        .Z(n11028) );
  HS65_LL_NAND4ABX3 U13110 ( .A(n13369), .B(n11029), .C(n11055), .D(n11028), 
        .Z(n11032) );
  HS65_LL_NAND4ABX3 U13111 ( .A(n11033), .B(n11032), .C(n11031), .D(n11030), 
        .Z(n11069) );
  HS65_LL_NAND3X2 U13112 ( .A(n11035), .B(n11034), .C(n13381), .Z(n11036) );
  HS65_LL_NOR4ABX2 U13113 ( .A(n11055), .B(n11037), .C(n11043), .D(n11036), 
        .Z(n11038) );
  HS65_LL_NAND3X2 U13114 ( .A(n11040), .B(n11039), .C(n11038), .Z(n11067) );
  HS65_LL_NAND4ABX3 U13115 ( .A(n11044), .B(n11043), .C(n11042), .D(n11041), 
        .Z(n11047) );
  HS65_LL_NAND4ABX3 U13116 ( .A(n11048), .B(n11047), .C(n11046), .D(n11045), 
        .Z(n13404) );
  HS65_LL_NOR4ABX2 U13117 ( .A(n11049), .B(n13384), .C(n13383), .D(n13404), 
        .Z(n11053) );
  HS65_LL_NOR4ABX2 U13118 ( .A(n11053), .B(n11052), .C(n11051), .D(n11050), 
        .Z(n11054) );
  HS65_LL_NAND3X2 U13119 ( .A(n11056), .B(n11055), .C(n11054), .Z(n11066) );
  HS65_LL_NAND4ABX3 U13120 ( .A(n11060), .B(n11059), .C(n11058), .D(n11057), 
        .Z(n11063) );
  HS65_LL_NOR2X2 U13121 ( .A(n13388), .B(n13387), .Z(n11061) );
  HS65_LL_NAND4ABX3 U13122 ( .A(n11064), .B(n11063), .C(n11062), .D(n11061), 
        .Z(n11065) );
  HS65_LL_MX41X4 U13123 ( .D0(n11069), .S0(n11068), .D1(n11067), .S1(n13393), 
        .D2(n11066), .S2(n13401), .D3(n11065), .S3(n13410), .Z(n15269) );
  HS65_LL_NOR4ABX2 U13124 ( .A(n11789), .B(n11071), .C(n11070), .D(n11577), 
        .Z(n11072) );
  HS65_LL_NAND3X2 U13125 ( .A(n11073), .B(n11072), .C(n11092), .Z(n14409) );
  HS65_LL_NOR2X2 U13126 ( .A(n11074), .B(n11798), .Z(n11076) );
  HS65_LL_NOR2X2 U13127 ( .A(n14438), .B(n14437), .Z(n11075) );
  HS65_LL_NAND4ABX3 U13128 ( .A(n11774), .B(n14409), .C(n11076), .D(n11075), 
        .Z(n11080) );
  HS65_LL_AOI12X2 U13129 ( .A(n11078), .B(n11077), .C(n11580), .Z(n11079) );
  HS65_LL_NAND4ABX3 U13130 ( .A(n11096), .B(n11080), .C(n11079), .D(n11802), 
        .Z(n11104) );
  HS65_LL_IVX2 U13131 ( .A(n11792), .Z(n11081) );
  HS65_LL_NOR2X2 U13132 ( .A(n11805), .B(n11081), .Z(n11599) );
  HS65_LL_NOR4ABX2 U13133 ( .A(n11083), .B(n11082), .C(n14446), .D(n11096), 
        .Z(n11084) );
  HS65_LL_NAND4ABX3 U13134 ( .A(n11086), .B(n11085), .C(n11599), .D(n11084), 
        .Z(n11103) );
  HS65_LL_IVX2 U13135 ( .A(n11611), .Z(n14451) );
  HS65_LL_NOR4ABX2 U13136 ( .A(n11565), .B(n11087), .C(n11597), .D(n11581), 
        .Z(n11088) );
  HS65_LL_NAND4ABX3 U13137 ( .A(n11572), .B(n14426), .C(n11089), .D(n11088), 
        .Z(n11102) );
  HS65_LL_AOI112X2 U13138 ( .A(n11091), .B(n11090), .C(n11577), .D(n11569), 
        .Z(n11098) );
  HS65_LL_IVX2 U13139 ( .A(n11573), .Z(n11093) );
  HS65_LL_NAND2X2 U13140 ( .A(n11093), .B(n11092), .Z(n14421) );
  HS65_LL_NAND4ABX3 U13141 ( .A(n11597), .B(n11096), .C(n11095), .D(n11094), 
        .Z(n11097) );
  HS65_LL_NOR4ABX2 U13142 ( .A(n11098), .B(n14419), .C(n14421), .D(n11097), 
        .Z(n11099) );
  HS65_LL_NAND3X2 U13143 ( .A(n14432), .B(n11100), .C(n11099), .Z(n11101) );
  HS65_LL_MX41X4 U13144 ( .D0(n11104), .S0(n14453), .D1(n11103), .S1(n14451), 
        .D2(n11102), .S2(n14449), .D3(n11101), .S3(n14447), .Z(n15129) );
  HS65_LL_MUXI21X2 U13145 ( .D0(w1[29]), .D1(n15128), .S0(n12148), .Z(n11105)
         );
  HS65_LLS_XOR3X2 U13146 ( .A(n15269), .B(n15129), .C(n11105), .Z(n11109) );
  HS65_LL_MUXI21X2 U13147 ( .D0(n15361), .D1(n14983), .S0(n15267), .Z(n14956)
         );
  HS65_LL_OAI21X2 U13148 ( .A(n14956), .B(n11109), .C(n14832), .Z(n11108) );
  HS65_LL_IVX2 U13149 ( .A(text_in_r[93]), .Z(n11106) );
  HS65_LL_OAI212X3 U13150 ( .A(w1[29]), .B(text_in_r[93]), .C(n15128), .D(
        n11106), .E(n15545), .Z(n11107) );
  HS65_LL_CBI4I1X3 U13151 ( .A(n11109), .B(n14956), .C(n11108), .D(n11107), 
        .Z(N215) );
  HS65_LL_IVX4 U13152 ( .A(n14808), .Z(n15727) );
  HS65_LL_OAI21X2 U13153 ( .A(w1[15]), .B(text_in_r[79]), .C(n15727), .Z(
        n11149) );
  HS65_LL_NAND2X2 U13154 ( .A(n11110), .B(n12178), .Z(n12840) );
  HS65_LL_NAND4ABX3 U13155 ( .A(n11124), .B(n12831), .C(n11112), .D(n11111), 
        .Z(n11114) );
  HS65_LL_NAND4ABX3 U13156 ( .A(n12840), .B(n11114), .C(n11113), .D(n14679), 
        .Z(n11144) );
  HS65_LL_AOI12X2 U13157 ( .A(n12168), .B(n11115), .C(n12183), .Z(n11121) );
  HS65_LL_NOR4ABX2 U13158 ( .A(n11119), .B(n11118), .C(n11117), .D(n11116), 
        .Z(n11120) );
  HS65_LL_NAND4ABX3 U13159 ( .A(n11123), .B(n11122), .C(n11121), .D(n11120), 
        .Z(n11143) );
  HS65_LL_NOR4ABX2 U13160 ( .A(n11126), .B(n12812), .C(n11125), .D(n11124), 
        .Z(n11134) );
  HS65_LL_NOR3X1 U13161 ( .A(n11129), .B(n11128), .C(n11127), .Z(n11132) );
  HS65_LL_NOR4ABX2 U13162 ( .A(n14650), .B(n11132), .C(n11131), .D(n11130), 
        .Z(n11133) );
  HS65_LL_NAND3X2 U13163 ( .A(n11135), .B(n11134), .C(n11133), .Z(n11142) );
  HS65_LL_NAND2X2 U13164 ( .A(n12154), .B(n12811), .Z(n11136) );
  HS65_LL_NOR3X1 U13165 ( .A(n12183), .B(n11137), .C(n11136), .Z(n11138) );
  HS65_LL_NAND4ABX3 U13166 ( .A(n11140), .B(n14664), .C(n11139), .D(n11138), 
        .Z(n11141) );
  HS65_LL_MX41X4 U13167 ( .D0(n11144), .S0(n12192), .D1(n11143), .S1(n14691), 
        .D2(n11142), .S2(n14683), .D3(n11141), .S3(n14685), .Z(n15443) );
  HS65_LL_IVX2 U13168 ( .A(n15443), .Z(n15444) );
  HS65_LL_IVX2 U13169 ( .A(w1[15]), .Z(n15014) );
  HS65_LL_MUXI21X2 U13170 ( .D0(w1[15]), .D1(n15014), .S0(n15445), .Z(n11145)
         );
  HS65_LL_MUXI21X2 U13171 ( .D0(n14955), .D1(n15359), .S0(n11145), .Z(n11146)
         );
  HS65_LL_MUXI21X2 U13172 ( .D0(n15443), .D1(n15444), .S0(n11146), .Z(n11147)
         );
  HS65_LL_MUXI21X2 U13173 ( .D0(n14843), .D1(n14842), .S0(n11147), .Z(n11148)
         );
  HS65_LL_CBI4I1X3 U13174 ( .A(text_in_r[79]), .B(w1[15]), .C(n11149), .D(
        n11148), .Z(N185) );
  HS65_LL_IVX4 U13175 ( .A(n14808), .Z(n15734) );
  HS65_LL_OAI21X2 U13176 ( .A(w0[15]), .B(text_in_r[111]), .C(n15734), .Z(
        n11353) );
  HS65_LL_OAI21X2 U13177 ( .A(n12554), .B(n12555), .C(n11171), .Z(n12866) );
  HS65_LL_NOR2X2 U13178 ( .A(n11187), .B(n11150), .Z(n14100) );
  HS65_LL_NOR2X2 U13179 ( .A(n14100), .B(n12546), .Z(n13466) );
  HS65_LL_NAND3AX3 U13180 ( .A(n12866), .B(n11151), .C(n13466), .Z(n14017) );
  HS65_LL_NOR2X2 U13181 ( .A(n12583), .B(n14001), .Z(n13480) );
  HS65_LL_NAND2X2 U13182 ( .A(n11152), .B(n12865), .Z(n13489) );
  HS65_LL_IVX2 U13183 ( .A(n11175), .Z(n13995) );
  HS65_LL_NAND2X2 U13184 ( .A(n13489), .B(n13995), .Z(n12886) );
  HS65_LL_NOR4ABX2 U13185 ( .A(n13480), .B(n13681), .C(n12549), .D(n12886), 
        .Z(n11153) );
  HS65_LL_NAND4ABX3 U13186 ( .A(n13474), .B(n14017), .C(n13994), .D(n11153), 
        .Z(n11194) );
  HS65_LL_NAND2AX4 U13187 ( .A(n12564), .B(n13489), .Z(n12577) );
  HS65_LL_OAI32X2 U13188 ( .A(n11156), .B(n13693), .C(n11183), .D(n11155), .E(
        n11154), .Z(n11157) );
  HS65_LL_OR3X4 U13189 ( .A(n13683), .B(n14096), .C(n11157), .Z(n11158) );
  HS65_LL_NAND4ABX3 U13190 ( .A(n14104), .B(n11158), .C(n12545), .D(n12894), 
        .Z(n11168) );
  HS65_LL_AOI12X2 U13191 ( .A(n11160), .B(n11159), .C(n14097), .Z(n11166) );
  HS65_LL_NOR3X1 U13192 ( .A(n13672), .B(n12582), .C(n14004), .Z(n14103) );
  HS65_LL_IVX2 U13193 ( .A(n12579), .Z(n12562) );
  HS65_LL_NOR2X2 U13194 ( .A(n11161), .B(n13677), .Z(n12543) );
  HS65_LL_IVX2 U13195 ( .A(n11162), .Z(n13990) );
  HS65_LL_NOR2X2 U13196 ( .A(n13990), .B(n11178), .Z(n12895) );
  HS65_LL_NAND2X2 U13197 ( .A(sa00[5]), .B(n11163), .Z(n14101) );
  HS65_LL_NAND2X2 U13198 ( .A(n13480), .B(n14101), .Z(n12879) );
  HS65_LL_NOR3X1 U13199 ( .A(n11164), .B(n12874), .C(n12879), .Z(n11165) );
  HS65_LL_NAND3X2 U13200 ( .A(n12543), .B(n12895), .C(n11165), .Z(n14018) );
  HS65_LL_NOR4ABX2 U13201 ( .A(n11166), .B(n14103), .C(n12562), .D(n14018), 
        .Z(n14106) );
  HS65_LL_NAND4ABX3 U13202 ( .A(n12577), .B(n11168), .C(n11167), .D(n14106), 
        .Z(n11193) );
  HS65_LL_NOR2X2 U13203 ( .A(n14108), .B(n11183), .Z(n14025) );
  HS65_LL_NOR2X2 U13204 ( .A(n13990), .B(n11169), .Z(n12890) );
  HS65_LL_IVX2 U13205 ( .A(n12548), .Z(n12880) );
  HS65_LL_NAND2X2 U13206 ( .A(n12880), .B(n13685), .Z(n12591) );
  HS65_LL_IVX2 U13207 ( .A(n12591), .Z(n14107) );
  HS65_LL_NOR4ABX2 U13208 ( .A(n11171), .B(n12588), .C(n11170), .D(n13683), 
        .Z(n11172) );
  HS65_LL_NAND3X2 U13209 ( .A(n12890), .B(n14107), .C(n11172), .Z(n14139) );
  HS65_LL_NAND2X2 U13210 ( .A(n11173), .B(n12884), .Z(n12892) );
  HS65_LL_NOR3X1 U13211 ( .A(n11175), .B(n11174), .C(n12892), .Z(n14111) );
  HS65_LL_NAND2X2 U13212 ( .A(n12894), .B(n14013), .Z(n12576) );
  HS65_LL_NOR2X2 U13213 ( .A(n11177), .B(n11176), .Z(n13472) );
  HS65_LL_NOR3X1 U13214 ( .A(n14096), .B(n13467), .C(n14012), .Z(n12581) );
  HS65_LL_NAND4ABX3 U13215 ( .A(n14097), .B(n11178), .C(n12581), .D(n14114), 
        .Z(n13686) );
  HS65_LL_NOR3X1 U13216 ( .A(n13472), .B(n13686), .C(n12879), .Z(n11179) );
  HS65_LL_OAI112X1 U13217 ( .A(n12554), .B(n11180), .C(n11179), .D(n13986), 
        .Z(n13492) );
  HS65_LL_NOR3X1 U13218 ( .A(n12576), .B(n13492), .C(n11181), .Z(n11182) );
  HS65_LL_NAND4ABX3 U13219 ( .A(n14025), .B(n14139), .C(n14111), .D(n11182), 
        .Z(n11192) );
  HS65_LL_OAI21X2 U13220 ( .A(n11184), .B(n11183), .C(n12560), .Z(n11186) );
  HS65_LL_NAND4ABX3 U13221 ( .A(n13478), .B(n11186), .C(n11185), .D(n13489), 
        .Z(n11189) );
  HS65_LL_NOR2X2 U13222 ( .A(n11188), .B(n11187), .Z(n13687) );
  HS65_LL_NOR2X2 U13223 ( .A(n12548), .B(n13687), .Z(n13669) );
  HS65_LL_NAND4ABX3 U13224 ( .A(n11190), .B(n11189), .C(n14111), .D(n13669), 
        .Z(n11191) );
  HS65_LL_MX41X4 U13225 ( .D0(n11194), .S0(n13709), .D1(n11193), .S1(n14130), 
        .D2(n11192), .S2(n14008), .D3(n11191), .S3(n14137), .Z(n15111) );
  HS65_LL_IVX2 U13226 ( .A(n15111), .Z(n15112) );
  HS65_LL_NAND3X2 U13227 ( .A(n12406), .B(n11195), .C(n11643), .Z(n11199) );
  HS65_LL_NOR4ABX2 U13228 ( .A(n11636), .B(n12954), .C(n13003), .D(n12997), 
        .Z(n11198) );
  HS65_LL_IVX2 U13229 ( .A(n12955), .Z(n13592) );
  HS65_LL_NOR3X1 U13230 ( .A(n12417), .B(n13592), .C(n11641), .Z(n13581) );
  HS65_LL_NOR4ABX2 U13231 ( .A(n13581), .B(n11203), .C(n12999), .D(n11196), 
        .Z(n11197) );
  HS65_LL_NAND4ABX3 U13232 ( .A(n11200), .B(n11199), .C(n11198), .D(n11197), 
        .Z(n11229) );
  HS65_LL_NAND2X2 U13233 ( .A(n11202), .B(n11201), .Z(n11648) );
  HS65_LL_OAI21X2 U13234 ( .A(n11649), .B(n11650), .C(n11203), .Z(n13589) );
  HS65_LL_NAND3X2 U13235 ( .A(n12418), .B(n13943), .C(n11204), .Z(n11205) );
  HS65_LL_NOR3X1 U13236 ( .A(n11206), .B(n13589), .C(n11205), .Z(n12427) );
  HS65_LL_OAI21X2 U13237 ( .A(n11208), .B(n11207), .C(n11631), .Z(n12972) );
  HS65_LL_NOR4ABX2 U13238 ( .A(n12427), .B(n11209), .C(n13942), .D(n12972), 
        .Z(n11210) );
  HS65_LL_OAI21X2 U13239 ( .A(n12986), .B(n12985), .C(n11210), .Z(n12968) );
  HS65_LL_NAND4ABX3 U13240 ( .A(n11211), .B(n12968), .C(n12959), .D(n13582), 
        .Z(n11213) );
  HS65_LL_NOR2X2 U13241 ( .A(n11625), .B(n13960), .Z(n13600) );
  HS65_LL_NAND4ABX3 U13242 ( .A(n11648), .B(n11213), .C(n11212), .D(n13600), 
        .Z(n11228) );
  HS65_LL_OAI13X1 U13243 ( .A(sa11[1]), .B(n11215), .C(n13578), .D(n11214), 
        .Z(n11218) );
  HS65_LL_NOR4ABX2 U13244 ( .A(n13582), .B(n13593), .C(n11625), .D(n11216), 
        .Z(n11217) );
  HS65_LL_NAND4ABX3 U13245 ( .A(n11219), .B(n11218), .C(n12401), .D(n11217), 
        .Z(n11227) );
  HS65_LL_AOI12X2 U13246 ( .A(n11221), .B(n11220), .C(n13605), .Z(n11627) );
  HS65_LL_IVX2 U13247 ( .A(n12398), .Z(n11222) );
  HS65_LL_NAND4ABX3 U13248 ( .A(n13598), .B(n11223), .C(n11627), .D(n11222), 
        .Z(n13954) );
  HS65_LL_NAND4ABX3 U13249 ( .A(n13612), .B(n11224), .C(n13610), .D(n11631), 
        .Z(n11225) );
  HS65_LL_NOR2X2 U13250 ( .A(n12962), .B(n11641), .Z(n12980) );
  HS65_LL_NAND4ABX3 U13251 ( .A(n13954), .B(n11225), .C(n12430), .D(n12980), 
        .Z(n11226) );
  HS65_LL_MX41X4 U13252 ( .D0(n11229), .S0(n13961), .D1(n11228), .S1(n13972), 
        .D2(n11227), .S2(n13614), .D3(n11226), .S3(n13981), .Z(n15251) );
  HS65_LL_MUXI21X2 U13253 ( .D0(n15112), .D1(n15111), .S0(n15251), .Z(n11230)
         );
  HS65_LL_NOR2X2 U13254 ( .A(n14822), .B(n11230), .Z(n14804) );
  HS65_LL_NOR2AX3 U13255 ( .A(n11230), .B(n15698), .Z(n14803) );
  HS65_LL_NAND2X2 U13256 ( .A(n11231), .B(n11240), .Z(n12622) );
  HS65_LL_NAND2X2 U13257 ( .A(n11708), .B(n12622), .Z(n14053) );
  HS65_LL_NOR2X2 U13258 ( .A(n13640), .B(n11276), .Z(n11724) );
  HS65_LL_NAND3X2 U13259 ( .A(n11724), .B(n11279), .C(n14031), .Z(n11232) );
  HS65_LL_NOR2X2 U13260 ( .A(n13558), .B(n11287), .Z(n11284) );
  HS65_LL_NOR2X2 U13261 ( .A(n11290), .B(n11284), .Z(n11277) );
  HS65_LL_NOR3X1 U13262 ( .A(n11278), .B(n11712), .C(n14054), .Z(n14064) );
  HS65_LL_NAND4ABX3 U13263 ( .A(n11285), .B(n11232), .C(n11277), .D(n14064), 
        .Z(n11233) );
  HS65_LL_NOR4ABX2 U13264 ( .A(n11234), .B(n11249), .C(n14053), .D(n11233), 
        .Z(n11265) );
  HS65_LL_IVX2 U13265 ( .A(n13657), .Z(n14071) );
  HS65_LL_AOI12X2 U13266 ( .A(n14058), .B(n11297), .C(n14039), .Z(n12632) );
  HS65_LL_NOR4ABX2 U13267 ( .A(n11235), .B(n13618), .C(n13541), .D(n12632), 
        .Z(n13644) );
  HS65_LL_NAND4ABX3 U13268 ( .A(n11252), .B(n11713), .C(n13644), .D(n11720), 
        .Z(n11236) );
  HS65_LL_AOI12X2 U13269 ( .A(n12625), .B(n12611), .C(n11236), .Z(n14073) );
  HS65_LL_NAND2X2 U13270 ( .A(n11237), .B(n11239), .Z(n12626) );
  HS65_LL_NAND2X2 U13271 ( .A(n13528), .B(n12626), .Z(n13646) );
  HS65_LL_NOR4ABX2 U13272 ( .A(n12615), .B(n14073), .C(n11712), .D(n13646), 
        .Z(n11238) );
  HS65_LL_NAND4ABX3 U13273 ( .A(n11291), .B(n12598), .C(n11238), .D(n13632), 
        .Z(n11255) );
  HS65_LL_NOR3X1 U13274 ( .A(n11285), .B(n14048), .C(n13529), .Z(n13634) );
  HS65_LL_NAND2X2 U13275 ( .A(n11240), .B(n11239), .Z(n14051) );
  HS65_LL_NAND4ABX3 U13276 ( .A(n11717), .B(n11241), .C(n13527), .D(n14051), 
        .Z(n11242) );
  HS65_LL_NOR3X1 U13277 ( .A(n13551), .B(n11284), .C(n11242), .Z(n11298) );
  HS65_LL_OAI21X2 U13278 ( .A(n11243), .B(n11293), .C(n12617), .Z(n11267) );
  HS65_LL_NOR3X1 U13279 ( .A(n14044), .B(n11244), .C(n11267), .Z(n11245) );
  HS65_LL_NAND4ABX3 U13280 ( .A(n11247), .B(n11246), .C(n11245), .D(n13641), 
        .Z(n13524) );
  HS65_LL_NOR2X2 U13281 ( .A(n11278), .B(n13524), .Z(n13547) );
  HS65_LL_NAND2AX4 U13282 ( .A(n13650), .B(n11727), .Z(n12597) );
  HS65_LL_NOR2X2 U13283 ( .A(n13533), .B(n12597), .Z(n13642) );
  HS65_LL_NAND2X2 U13284 ( .A(n11248), .B(n12626), .Z(n11273) );
  HS65_LL_NOR3X1 U13285 ( .A(n11712), .B(n13515), .C(n11273), .Z(n11250) );
  HS65_LL_NAND3X2 U13286 ( .A(n11251), .B(n11250), .C(n11249), .Z(n12603) );
  HS65_LL_NOR4ABX2 U13287 ( .A(n13547), .B(n13642), .C(n11252), .D(n12603), 
        .Z(n11253) );
  HS65_LL_AOI13X2 U13288 ( .A(n13634), .B(n11298), .C(n11253), .D(n14079), .Z(
        n11254) );
  HS65_LL_CBI4I6X2 U13289 ( .A(n11256), .B(n11255), .C(n14067), .D(n11254), 
        .Z(n11264) );
  HS65_LL_NOR2X2 U13290 ( .A(n13629), .B(n13646), .Z(n11300) );
  HS65_LL_NOR4ABX2 U13291 ( .A(n13544), .B(n14028), .C(n13630), .D(n13526), 
        .Z(n11257) );
  HS65_LL_NAND4ABX3 U13292 ( .A(n13650), .B(n12606), .C(n11300), .D(n11257), 
        .Z(n11731) );
  HS65_LL_OAI21X2 U13293 ( .A(n11721), .B(n11258), .C(n11714), .Z(n12624) );
  HS65_LL_NAND4ABX3 U13294 ( .A(n11290), .B(n12624), .C(n11259), .D(n13626), 
        .Z(n11706) );
  HS65_LL_OAI112X1 U13295 ( .A(sa33[1]), .B(n14031), .C(n11260), .D(n12615), 
        .Z(n11261) );
  HS65_LL_NAND4ABX3 U13296 ( .A(n11267), .B(n11261), .C(n13621), .D(n11702), 
        .Z(n11262) );
  HS65_LL_OAI13X1 U13297 ( .A(n11731), .B(n11706), .C(n11262), .D(n14075), .Z(
        n11263) );
  HS65_LL_OAI112X1 U13298 ( .A(n11265), .B(n14071), .C(n11264), .D(n11263), 
        .Z(n15435) );
  HS65_LL_IVX2 U13299 ( .A(n15435), .Z(n15436) );
  HS65_LL_NOR2X2 U13300 ( .A(n12629), .B(n12597), .Z(n13512) );
  HS65_LL_AOI12X2 U13301 ( .A(n13517), .B(n13518), .C(n13533), .Z(n11711) );
  HS65_LL_NOR3AX2 U13302 ( .A(sa33[7]), .B(n11266), .C(n13558), .Z(n11269) );
  HS65_LL_OAI21X2 U13303 ( .A(n11721), .B(n11293), .C(n11702), .Z(n13540) );
  HS65_LL_NAND4ABX3 U13304 ( .A(n11267), .B(n13540), .C(n13548), .D(n12600), 
        .Z(n11268) );
  HS65_LL_NOR4ABX2 U13305 ( .A(n14064), .B(n13528), .C(n11269), .D(n11268), 
        .Z(n12604) );
  HS65_LL_NOR2X2 U13306 ( .A(n14044), .B(n13537), .Z(n13620) );
  HS65_LL_NAND2X2 U13307 ( .A(n11275), .B(n11270), .Z(n14041) );
  HS65_LL_NOR4ABX2 U13308 ( .A(n13527), .B(n14041), .C(n11291), .D(n11290), 
        .Z(n11271) );
  HS65_LL_NAND3X2 U13309 ( .A(n11272), .B(n11271), .C(n11289), .Z(n11719) );
  HS65_LL_NOR4ABX2 U13310 ( .A(n12604), .B(n13620), .C(n11273), .D(n11719), 
        .Z(n11274) );
  HS65_LL_NAND3X2 U13311 ( .A(n13512), .B(n11711), .C(n11274), .Z(n11306) );
  HS65_LL_IVX2 U13312 ( .A(n14079), .Z(n13659) );
  HS65_LL_AOI12X2 U13313 ( .A(n14036), .B(n11275), .C(n13630), .Z(n11704) );
  HS65_LL_IVX2 U13314 ( .A(n11276), .Z(n11707) );
  HS65_LL_NAND3AX3 U13315 ( .A(n13526), .B(n11277), .C(n11707), .Z(n12616) );
  HS65_LL_NOR4ABX2 U13316 ( .A(n11704), .B(n11279), .C(n11278), .D(n12616), 
        .Z(n11280) );
  HS65_LL_NAND3X2 U13317 ( .A(n11281), .B(n14073), .C(n11280), .Z(n13550) );
  HS65_LL_IVX2 U13318 ( .A(n12606), .Z(n12620) );
  HS65_LL_NOR4ABX2 U13319 ( .A(n12620), .B(n12626), .C(n11712), .D(n14034), 
        .Z(n14056) );
  HS65_LL_NAND4ABX3 U13320 ( .A(n11283), .B(n13550), .C(n11282), .D(n14056), 
        .Z(n11305) );
  HS65_LL_IVX2 U13321 ( .A(n11284), .Z(n13539) );
  HS65_LL_NOR2X2 U13322 ( .A(n11285), .B(n13529), .Z(n11286) );
  HS65_LL_NAND4ABX3 U13323 ( .A(n13551), .B(n14044), .C(n13539), .D(n11286), 
        .Z(n11730) );
  HS65_LL_NOR2X2 U13324 ( .A(n11287), .B(n11725), .Z(n13553) );
  HS65_LL_NOR2X2 U13325 ( .A(n11288), .B(n13553), .Z(n13538) );
  HS65_LL_NAND4ABX3 U13326 ( .A(n13543), .B(n13526), .C(n13538), .D(n11289), 
        .Z(n11296) );
  HS65_LL_NOR2X2 U13327 ( .A(n11291), .B(n11290), .Z(n11294) );
  HS65_LL_OAI112X1 U13328 ( .A(n11293), .B(n14039), .C(n11292), .D(n14041), 
        .Z(n13649) );
  HS65_LL_NOR4ABX2 U13329 ( .A(n11300), .B(n11294), .C(n14054), .D(n13649), 
        .Z(n11295) );
  HS65_LL_NAND3X2 U13330 ( .A(n11295), .B(n11702), .C(n12622), .Z(n13624) );
  HS65_LL_NOR3X1 U13331 ( .A(n12629), .B(n12597), .C(n13624), .Z(n11709) );
  HS65_LL_NAND4ABX3 U13332 ( .A(n11730), .B(n11296), .C(n11301), .D(n11709), 
        .Z(n11304) );
  HS65_LL_NAND2X2 U13333 ( .A(n12612), .B(n13544), .Z(n12630) );
  HS65_LL_OAI21X2 U13334 ( .A(n14039), .B(n11297), .C(n13632), .Z(n14033) );
  HS65_LL_NAND2X2 U13335 ( .A(n13548), .B(n12600), .Z(n11299) );
  HS65_LL_NAND4ABX3 U13336 ( .A(n14033), .B(n11299), .C(n13654), .D(n11298), 
        .Z(n11302) );
  HS65_LL_NAND4ABX3 U13337 ( .A(n12630), .B(n11302), .C(n11301), .D(n11300), 
        .Z(n11303) );
  HS65_LL_MX41X4 U13338 ( .D0(n11306), .S0(n13659), .D1(n11305), .S1(n13657), 
        .D2(n11304), .S2(n14067), .D3(n11303), .S3(n14075), .Z(n15531) );
  HS65_LL_IVX2 U13339 ( .A(n15531), .Z(n15530) );
  HS65_LL_NOR2X2 U13340 ( .A(n12485), .B(n11307), .Z(n12480) );
  HS65_LL_NOR2X2 U13341 ( .A(n11308), .B(n11756), .Z(n11320) );
  HS65_LL_NAND3X2 U13342 ( .A(n12480), .B(n11320), .C(n12458), .Z(n11750) );
  HS65_LL_NAND2X2 U13343 ( .A(n11309), .B(n11340), .Z(n12447) );
  HS65_LL_IVX2 U13344 ( .A(n12447), .Z(n12536) );
  HS65_LL_OR2X4 U13345 ( .A(n11310), .B(n12453), .Z(n11671) );
  HS65_LL_NAND3X2 U13346 ( .A(sa22[5]), .B(sa22[0]), .C(n11311), .Z(n12450) );
  HS65_LL_NAND4ABX3 U13347 ( .A(n11671), .B(n12927), .C(n12450), .D(n12516), 
        .Z(n11312) );
  HS65_LL_NOR3X1 U13348 ( .A(n12536), .B(n12439), .C(n11312), .Z(n11314) );
  HS65_LL_NAND3X2 U13349 ( .A(n11314), .B(n11313), .C(n12506), .Z(n11760) );
  HS65_LL_NAND4ABX3 U13350 ( .A(n11325), .B(n11760), .C(n12454), .D(n12501), 
        .Z(n11317) );
  HS65_LL_NOR2X2 U13351 ( .A(n12530), .B(n12524), .Z(n11315) );
  HS65_LL_NAND4ABX3 U13352 ( .A(n11750), .B(n11317), .C(n11316), .D(n11315), 
        .Z(n11347) );
  HS65_LL_NOR4ABX2 U13353 ( .A(n11320), .B(n11319), .C(n11318), .D(n12469), 
        .Z(n11686) );
  HS65_LL_NOR4ABX2 U13354 ( .A(n11686), .B(n11331), .C(n12503), .D(n12907), 
        .Z(n11327) );
  HS65_LL_NOR2X2 U13355 ( .A(n11321), .B(n11751), .Z(n12478) );
  HS65_LL_OAI21X2 U13356 ( .A(n11324), .B(n11323), .C(n11322), .Z(n12510) );
  HS65_LL_NOR4ABX2 U13357 ( .A(n12478), .B(n12515), .C(n11325), .D(n12510), 
        .Z(n11326) );
  HS65_LL_NAND3X2 U13358 ( .A(n12457), .B(n11327), .C(n11326), .Z(n11346) );
  HS65_LL_NAND2X2 U13359 ( .A(n12533), .B(n12458), .Z(n11338) );
  HS65_LL_NOR3X1 U13360 ( .A(n11343), .B(n12524), .C(n11328), .Z(n11329) );
  HS65_LL_NAND3X2 U13361 ( .A(n11690), .B(n11329), .C(n12447), .Z(n11742) );
  HS65_LL_NAND2AX4 U13362 ( .A(n12460), .B(n12506), .Z(n12928) );
  HS65_LL_NOR3X1 U13363 ( .A(n12446), .B(n12440), .C(n12928), .Z(n11694) );
  HS65_LL_NOR4ABX2 U13364 ( .A(n11694), .B(n11331), .C(n11743), .D(n11330), 
        .Z(n11332) );
  HS65_LL_NAND4ABX3 U13365 ( .A(n12504), .B(n11333), .C(n11332), .D(n12515), 
        .Z(n12471) );
  HS65_LL_NOR2X2 U13366 ( .A(n11334), .B(n12503), .Z(n11682) );
  HS65_LL_NOR3X1 U13367 ( .A(n11335), .B(n12530), .C(n12498), .Z(n12443) );
  HS65_LL_NAND3X2 U13368 ( .A(n11682), .B(n12443), .C(n12501), .Z(n11336) );
  HS65_LL_NOR3X1 U13369 ( .A(n11742), .B(n12471), .C(n11336), .Z(n11337) );
  HS65_LL_NAND4ABX3 U13370 ( .A(n12937), .B(n11338), .C(n11337), .D(n12531), 
        .Z(n11345) );
  HS65_LL_IVX2 U13371 ( .A(n11339), .Z(n12943) );
  HS65_LL_NAND2X2 U13372 ( .A(n12448), .B(n12473), .Z(n12921) );
  HS65_LL_AOI12X2 U13373 ( .A(n11340), .B(n12499), .C(n12921), .Z(n11341) );
  HS65_LL_NAND4ABX3 U13374 ( .A(n11343), .B(n12503), .C(n11342), .D(n11341), 
        .Z(n11344) );
  HS65_LL_MX41X4 U13375 ( .D0(n11347), .S0(n12540), .D1(n11346), .S1(n12951), 
        .D2(n11345), .S2(n12943), .D3(n11344), .S3(n12945), .Z(n15347) );
  HS65_LL_MUXI21X2 U13376 ( .D0(w0[15]), .D1(n11348), .S0(n15347), .Z(n11349)
         );
  HS65_LL_MUXI21X2 U13377 ( .D0(n15531), .D1(n15530), .S0(n11349), .Z(n11350)
         );
  HS65_LL_MUXI21X2 U13378 ( .D0(n15435), .D1(n15436), .S0(n11350), .Z(n11351)
         );
  HS65_LL_MUXI21X2 U13379 ( .D0(n14804), .D1(n14803), .S0(n11351), .Z(n11352)
         );
  HS65_LL_CBI4I1X3 U13380 ( .A(text_in_r[111]), .B(w0[15]), .C(n11353), .D(
        n11352), .Z(N249) );
  HS65_LL_IVX2 U13381 ( .A(sa21[7]), .Z(n11369) );
  HS65_LL_NAND2X2 U13382 ( .A(sa21[1]), .B(n11369), .Z(n11354) );
  HS65_LL_IVX2 U13383 ( .A(sa21[5]), .Z(n11359) );
  HS65_LL_NAND3X2 U13384 ( .A(sa21[0]), .B(sa21[3]), .C(n11359), .Z(n11363) );
  HS65_LL_NOR2X2 U13385 ( .A(n11354), .B(n11363), .Z(n11915) );
  HS65_LL_IVX2 U13386 ( .A(sa21[0]), .Z(n11358) );
  HS65_LL_NOR2X2 U13387 ( .A(sa21[3]), .B(n11358), .Z(n11911) );
  HS65_LL_NOR3X1 U13388 ( .A(sa21[6]), .B(sa21[1]), .C(n11369), .Z(n12677) );
  HS65_LL_NAND3X2 U13389 ( .A(sa21[5]), .B(n11911), .C(n12677), .Z(n13220) );
  HS65_LL_IVX2 U13390 ( .A(sa21[6]), .Z(n13826) );
  HS65_LL_NOR2X2 U13391 ( .A(n13826), .B(n11354), .Z(n12644) );
  HS65_LL_NAND2X2 U13392 ( .A(sa21[3]), .B(n11358), .Z(n12642) );
  HS65_LL_NOR2X2 U13393 ( .A(n11359), .B(n12642), .Z(n11923) );
  HS65_LL_NAND2X2 U13394 ( .A(n12644), .B(n11923), .Z(n11938) );
  HS65_LL_NAND2X2 U13395 ( .A(n13220), .B(n11938), .Z(n13838) );
  HS65_LL_NOR2X2 U13396 ( .A(n11915), .B(n13838), .Z(n14271) );
  HS65_LL_NOR3X1 U13397 ( .A(sa21[1]), .B(n11369), .C(n13826), .Z(n11926) );
  HS65_LL_NAND2X2 U13398 ( .A(sa21[0]), .B(sa21[3]), .Z(n12674) );
  HS65_LL_NOR2X2 U13399 ( .A(n11359), .B(n12674), .Z(n11370) );
  HS65_LL_NAND2X2 U13400 ( .A(n11926), .B(n11370), .Z(n13210) );
  HS65_LL_NAND2X2 U13401 ( .A(n14271), .B(n13210), .Z(n13881) );
  HS65_LL_IVX2 U13402 ( .A(sa21[1]), .Z(n13825) );
  HS65_LL_NOR2X2 U13403 ( .A(sa21[5]), .B(n12642), .Z(n12659) );
  HS65_LL_IVX2 U13404 ( .A(n12659), .Z(n11382) );
  HS65_LL_NOR3X1 U13405 ( .A(n13825), .B(n11382), .C(sa21[6]), .Z(n11376) );
  HS65_LL_NAND2X2 U13406 ( .A(n12659), .B(n12644), .Z(n14247) );
  HS65_LL_NAND2X2 U13407 ( .A(n12677), .B(n11923), .Z(n14252) );
  HS65_LL_NAND2X2 U13408 ( .A(n14247), .B(n14252), .Z(n11924) );
  HS65_LL_NOR2X2 U13409 ( .A(sa21[0]), .B(sa21[3]), .Z(n11355) );
  HS65_LL_NAND2X2 U13410 ( .A(sa21[5]), .B(n11355), .Z(n11388) );
  HS65_LL_IVX2 U13411 ( .A(n11388), .Z(n11381) );
  HS65_LL_NOR2X2 U13412 ( .A(sa21[6]), .B(sa21[1]), .Z(n14152) );
  HS65_LL_NAND2X2 U13413 ( .A(n14152), .B(n11369), .Z(n11368) );
  HS65_LL_IVX2 U13414 ( .A(n11368), .Z(n11910) );
  HS65_LL_NAND2X2 U13415 ( .A(n11381), .B(n11910), .Z(n14240) );
  HS65_LL_NOR2X2 U13416 ( .A(sa21[6]), .B(n11354), .Z(n11384) );
  HS65_LL_NAND2X2 U13417 ( .A(n11355), .B(n11384), .Z(n14170) );
  HS65_LL_NAND4ABX3 U13418 ( .A(n11376), .B(n11924), .C(n14240), .D(n14170), 
        .Z(n11361) );
  HS65_LL_NAND3X2 U13419 ( .A(sa21[6]), .B(n11369), .C(n13825), .Z(n12675) );
  HS65_LL_NAND2X2 U13420 ( .A(n11911), .B(n11359), .Z(n13829) );
  HS65_LL_NOR2X2 U13421 ( .A(n12675), .B(n13829), .Z(n13233) );
  HS65_LL_NAND2X2 U13422 ( .A(n11355), .B(n11359), .Z(n11357) );
  HS65_LL_NAND3X2 U13423 ( .A(sa21[7]), .B(sa21[1]), .C(n13826), .Z(n11922) );
  HS65_LL_NOR2X2 U13424 ( .A(n11357), .B(n11922), .Z(n13879) );
  HS65_LL_NAND2X2 U13425 ( .A(sa21[5]), .B(n11911), .Z(n11942) );
  HS65_LL_NOR2X2 U13426 ( .A(n12675), .B(n11942), .Z(n13861) );
  HS65_LL_NAND3X2 U13427 ( .A(sa21[6]), .B(sa21[7]), .C(sa21[1]), .Z(n11941)
         );
  HS65_LL_IVX2 U13428 ( .A(n11923), .Z(n11373) );
  HS65_LL_NOR2X2 U13429 ( .A(n11941), .B(n11373), .Z(n11921) );
  HS65_LL_NOR2X2 U13430 ( .A(n13861), .B(n11921), .Z(n12661) );
  HS65_LL_IVX2 U13431 ( .A(n11942), .Z(n11371) );
  HS65_LL_NAND2X2 U13432 ( .A(n11371), .B(n12644), .Z(n11945) );
  HS65_LL_IVX2 U13433 ( .A(n11945), .Z(n12683) );
  HS65_LL_NAND2X2 U13434 ( .A(n11370), .B(n12644), .Z(n13206) );
  HS65_LL_IVX2 U13435 ( .A(n13829), .Z(n11380) );
  HS65_LL_NAND2X2 U13436 ( .A(n11380), .B(n11384), .Z(n12647) );
  HS65_LL_NAND2X2 U13437 ( .A(n13206), .B(n12647), .Z(n11913) );
  HS65_LL_NOR2X2 U13438 ( .A(n12683), .B(n11913), .Z(n14258) );
  HS65_LL_NOR2X2 U13439 ( .A(n11941), .B(n11363), .Z(n11374) );
  HS65_LL_IVX2 U13440 ( .A(n11926), .Z(n11387) );
  HS65_LL_NOR2X2 U13441 ( .A(n11387), .B(n11373), .Z(n14256) );
  HS65_LL_NOR2X2 U13442 ( .A(n11374), .B(n14256), .Z(n13806) );
  HS65_LL_NAND3X2 U13443 ( .A(n12661), .B(n14258), .C(n13806), .Z(n11356) );
  HS65_LL_NOR3X1 U13444 ( .A(n13233), .B(n13879), .C(n11356), .Z(n14272) );
  HS65_LL_NOR2X2 U13445 ( .A(n11388), .B(n11922), .Z(n13234) );
  HS65_LL_NOR2X2 U13446 ( .A(n13829), .B(n11941), .Z(n13867) );
  HS65_LL_IVX2 U13447 ( .A(n11357), .Z(n11385) );
  HS65_LL_NAND2X2 U13448 ( .A(n11910), .B(n11385), .Z(n13228) );
  HS65_LL_IVX2 U13449 ( .A(n12675), .Z(n14266) );
  HS65_LL_IVX2 U13450 ( .A(n11363), .Z(n14151) );
  HS65_LL_NAND2X2 U13451 ( .A(n14266), .B(n14151), .Z(n13235) );
  HS65_LL_NAND2X2 U13452 ( .A(n13228), .B(n13235), .Z(n14265) );
  HS65_LL_NOR2X2 U13453 ( .A(n13867), .B(n14265), .Z(n11362) );
  HS65_LL_NAND3X2 U13454 ( .A(sa21[0]), .B(sa21[3]), .C(n12677), .Z(n12652) );
  HS65_LL_NOR2X2 U13455 ( .A(n11387), .B(n11357), .Z(n13820) );
  HS65_LL_NAND3X2 U13456 ( .A(sa21[1]), .B(n11371), .C(n13826), .Z(n13214) );
  HS65_LL_IVX2 U13457 ( .A(n11922), .Z(n11365) );
  HS65_LL_NAND2X2 U13458 ( .A(n11370), .B(n11365), .Z(n11907) );
  HS65_LL_NAND2X2 U13459 ( .A(n14266), .B(n12659), .Z(n13876) );
  HS65_LL_NAND3X2 U13460 ( .A(n13214), .B(n11907), .C(n13876), .Z(n13871) );
  HS65_LL_NOR4ABX2 U13461 ( .A(n11362), .B(n12652), .C(n13820), .D(n13871), 
        .Z(n11360) );
  HS65_LL_NAND2X2 U13462 ( .A(n11380), .B(n12644), .Z(n13236) );
  HS65_LL_NAND3AX3 U13463 ( .A(sa21[3]), .B(n11358), .C(n12644), .Z(n11937) );
  HS65_LL_NOR2X2 U13464 ( .A(n11359), .B(n11937), .Z(n14154) );
  HS65_LL_IVX2 U13465 ( .A(n14154), .Z(n14238) );
  HS65_LL_NAND3X2 U13466 ( .A(n11360), .B(n13236), .C(n14238), .Z(n13223) );
  HS65_LL_NOR2X2 U13467 ( .A(n13234), .B(n13223), .Z(n13889) );
  HS65_LL_NAND4ABX3 U13468 ( .A(n13881), .B(n11361), .C(n14272), .D(n13889), 
        .Z(n11395) );
  HS65_LL_NOR2X2 U13469 ( .A(sa21[2]), .B(sa21[4]), .Z(n14285) );
  HS65_LL_IVX2 U13470 ( .A(n11370), .Z(n11379) );
  HS65_LL_NOR2X2 U13471 ( .A(n11379), .B(n11941), .Z(n13839) );
  HS65_LL_NOR2X2 U13472 ( .A(n11941), .B(n11382), .Z(n12689) );
  HS65_LL_IVX2 U13473 ( .A(n11938), .Z(n11383) );
  HS65_LL_NOR2X2 U13474 ( .A(n12689), .B(n11383), .Z(n14174) );
  HS65_LL_NAND2X2 U13475 ( .A(n12659), .B(n11384), .Z(n11375) );
  HS65_LL_NAND2X2 U13476 ( .A(n14174), .B(n11375), .Z(n13870) );
  HS65_LL_NAND2X2 U13477 ( .A(n11381), .B(n11384), .Z(n13818) );
  HS65_LL_AND2X4 U13478 ( .A(n13818), .B(n11362), .Z(n13218) );
  HS65_LL_NAND2X2 U13479 ( .A(n11926), .B(n11380), .Z(n12650) );
  HS65_LL_NAND4ABX3 U13480 ( .A(n13839), .B(n13870), .C(n13218), .D(n12650), 
        .Z(n14255) );
  HS65_LL_NAND2X2 U13481 ( .A(n11926), .B(n12659), .Z(n12680) );
  HS65_LL_NAND2X2 U13482 ( .A(n11380), .B(n11365), .Z(n13817) );
  HS65_LL_NAND2X2 U13483 ( .A(n12680), .B(n13817), .Z(n13866) );
  HS65_LL_NOR2X2 U13484 ( .A(n11388), .B(n12675), .Z(n14164) );
  HS65_LL_NAND2X2 U13485 ( .A(n11910), .B(n14151), .Z(n12651) );
  HS65_LL_NAND2AX4 U13486 ( .A(n14164), .B(n12651), .Z(n13215) );
  HS65_LL_NOR2X2 U13487 ( .A(n13866), .B(n13215), .Z(n14276) );
  HS65_LL_IVX2 U13488 ( .A(n13233), .Z(n12646) );
  HS65_LL_NAND2X2 U13489 ( .A(n14276), .B(n12646), .Z(n13222) );
  HS65_LL_NAND2X2 U13490 ( .A(n12677), .B(n11385), .Z(n11936) );
  HS65_LL_IVX2 U13491 ( .A(n11936), .Z(n13204) );
  HS65_LL_NOR2X2 U13492 ( .A(n13204), .B(n14256), .Z(n14244) );
  HS65_LL_NAND2X2 U13493 ( .A(n11384), .B(n11385), .Z(n13231) );
  HS65_LL_NAND2X2 U13494 ( .A(n14244), .B(n13231), .Z(n12649) );
  HS65_LL_NAND2X2 U13495 ( .A(n11371), .B(n11910), .Z(n12684) );
  HS65_LL_NAND2X2 U13496 ( .A(n14266), .B(n11385), .Z(n13828) );
  HS65_LL_NAND2X2 U13497 ( .A(n12684), .B(n13828), .Z(n14169) );
  HS65_LL_NAND2X2 U13498 ( .A(n11910), .B(n12659), .Z(n14257) );
  HS65_LL_NAND2X2 U13499 ( .A(n11380), .B(n11910), .Z(n13237) );
  HS65_LL_NAND2X2 U13500 ( .A(n14257), .B(n13237), .Z(n11932) );
  HS65_LL_NOR3X1 U13501 ( .A(n12649), .B(n14169), .C(n11932), .Z(n11364) );
  HS65_LL_NOR2X2 U13502 ( .A(sa21[5]), .B(n11937), .Z(n14177) );
  HS65_LL_AOI12X2 U13503 ( .A(n11388), .B(n11363), .C(n11941), .Z(n13878) );
  HS65_LL_NOR4ABX2 U13504 ( .A(n11364), .B(n14247), .C(n14177), .D(n13878), 
        .Z(n13874) );
  HS65_LL_NAND2X2 U13505 ( .A(n11911), .B(n12677), .Z(n11366) );
  HS65_LL_NAND2X2 U13506 ( .A(n14151), .B(n11365), .Z(n13209) );
  HS65_LL_AND2X4 U13507 ( .A(n11384), .B(n14151), .Z(n14270) );
  HS65_LL_NAND2X2 U13508 ( .A(n14240), .B(n14238), .Z(n11931) );
  HS65_LL_NOR4ABX2 U13509 ( .A(n11366), .B(n13209), .C(n14270), .D(n11931), 
        .Z(n11367) );
  HS65_LL_NAND4ABX3 U13510 ( .A(n14255), .B(n13222), .C(n13874), .D(n11367), 
        .Z(n11394) );
  HS65_LL_IVX2 U13511 ( .A(sa21[2]), .Z(n11391) );
  HS65_LL_NOR2X2 U13512 ( .A(sa21[4]), .B(n11391), .Z(n14283) );
  HS65_LL_NAND2X2 U13513 ( .A(n11370), .B(n11384), .Z(n13221) );
  HS65_LL_IVX2 U13514 ( .A(n13221), .Z(n13845) );
  HS65_LL_NAND2X2 U13515 ( .A(n12677), .B(n12659), .Z(n12648) );
  HS65_LL_NOR2X2 U13516 ( .A(n11368), .B(n12642), .Z(n13213) );
  HS65_LL_NAND2X2 U13517 ( .A(sa21[5]), .B(n13213), .Z(n12670) );
  HS65_LL_NAND2X2 U13518 ( .A(n12648), .B(n12670), .Z(n12663) );
  HS65_LL_NAND3X2 U13519 ( .A(sa21[6]), .B(n12659), .C(n11369), .Z(n11935) );
  HS65_LL_NAND4ABX3 U13520 ( .A(n13845), .B(n12663), .C(n11935), .D(n12652), 
        .Z(n13242) );
  HS65_LL_IVX2 U13521 ( .A(n13861), .Z(n12656) );
  HS65_LL_NAND2X2 U13522 ( .A(n11370), .B(n11910), .Z(n12664) );
  HS65_LL_NAND2X2 U13523 ( .A(n12656), .B(n12664), .Z(n12679) );
  HS65_LL_NAND2X2 U13524 ( .A(n11381), .B(n12677), .Z(n14166) );
  HS65_LL_NAND2X2 U13525 ( .A(n14266), .B(n11370), .Z(n11927) );
  HS65_LL_NAND2X2 U13526 ( .A(n14166), .B(n11927), .Z(n13891) );
  HS65_LL_NOR4ABX2 U13527 ( .A(n11945), .B(n13237), .C(n12679), .D(n13891), 
        .Z(n14178) );
  HS65_LL_IVX2 U13528 ( .A(n11907), .Z(n13211) );
  HS65_LL_NOR3X1 U13529 ( .A(n13234), .B(n14270), .C(n13211), .Z(n11934) );
  HS65_LL_NAND2X2 U13530 ( .A(n11371), .B(n11384), .Z(n11378) );
  HS65_LL_NOR4ABX2 U13531 ( .A(n11934), .B(n11378), .C(n13879), .D(n14169), 
        .Z(n11372) );
  HS65_LL_NAND4ABX3 U13532 ( .A(n14255), .B(n13242), .C(n14178), .D(n11372), 
        .Z(n11393) );
  HS65_LL_IVX2 U13533 ( .A(sa21[4]), .Z(n11390) );
  HS65_LL_NOR2X2 U13534 ( .A(sa21[2]), .B(n11390), .Z(n14281) );
  HS65_LL_NOR2X2 U13535 ( .A(n11922), .B(n11373), .Z(n13860) );
  HS65_LL_NOR2X2 U13536 ( .A(n13860), .B(n11374), .Z(n13887) );
  HS65_LL_NOR2X2 U13537 ( .A(sa21[5]), .B(n12652), .Z(n13835) );
  HS65_LL_NOR2X2 U13538 ( .A(n13835), .B(n13867), .Z(n11914) );
  HS65_LL_IVX2 U13539 ( .A(n11375), .Z(n14144) );
  HS65_LL_NAND2X2 U13540 ( .A(sa21[7]), .B(n11376), .Z(n14173) );
  HS65_LL_NAND2X2 U13541 ( .A(n13206), .B(n14173), .Z(n13875) );
  HS65_LL_NOR3X1 U13542 ( .A(n13204), .B(n14144), .C(n13875), .Z(n11377) );
  HS65_LL_NAND3X2 U13543 ( .A(n13887), .B(n11914), .C(n11377), .Z(n12668) );
  HS65_LL_IVX2 U13544 ( .A(n11378), .Z(n13840) );
  HS65_LL_NOR3X1 U13545 ( .A(sa21[6]), .B(sa21[1]), .C(n11379), .Z(n13200) );
  HS65_LL_NAND2X2 U13546 ( .A(n14151), .B(n12644), .Z(n13824) );
  HS65_LL_NOR2X2 U13547 ( .A(n11387), .B(n11942), .Z(n13239) );
  HS65_LL_NAND2X2 U13548 ( .A(n11380), .B(n12677), .Z(n14157) );
  HS65_LL_IVX2 U13549 ( .A(n11941), .Z(n11386) );
  HS65_LL_NAND2X2 U13550 ( .A(n11381), .B(n11386), .Z(n14239) );
  HS65_LL_NAND2X2 U13551 ( .A(n14157), .B(n14239), .Z(n12643) );
  HS65_LL_NOR2X2 U13552 ( .A(n13239), .B(n12643), .Z(n14167) );
  HS65_LL_NAND4ABX3 U13553 ( .A(n13840), .B(n13200), .C(n13824), .D(n14167), 
        .Z(n14261) );
  HS65_LL_NAND2X2 U13554 ( .A(n13231), .B(n12670), .Z(n13812) );
  HS65_LL_NOR4ABX2 U13555 ( .A(n12650), .B(n13236), .C(n11921), .D(n13812), 
        .Z(n14175) );
  HS65_LL_NOR3X1 U13556 ( .A(sa21[1]), .B(n13826), .C(n11382), .Z(n11928) );
  HS65_LL_NOR2X2 U13557 ( .A(n13839), .B(n11928), .Z(n13202) );
  HS65_LL_NOR2X2 U13558 ( .A(n13234), .B(n11383), .Z(n13833) );
  HS65_LL_NAND3X2 U13559 ( .A(sa21[5]), .B(sa21[3]), .C(n11384), .Z(n11940) );
  HS65_LL_NOR2X2 U13560 ( .A(sa21[0]), .B(n11940), .Z(n14246) );
  HS65_LL_NAND3X2 U13561 ( .A(n12648), .B(n11927), .C(n13228), .Z(n13207) );
  HS65_LL_NAND2X2 U13562 ( .A(n11386), .B(n11385), .Z(n13229) );
  HS65_LL_IVX2 U13563 ( .A(n12684), .Z(n13809) );
  HS65_LL_NOR2AX3 U13564 ( .A(n13229), .B(n13809), .Z(n12666) );
  HS65_LL_NOR2X2 U13565 ( .A(n11388), .B(n11387), .Z(n11943) );
  HS65_LL_NOR2AX3 U13566 ( .A(n13209), .B(n11943), .Z(n14179) );
  HS65_LL_NAND4ABX3 U13567 ( .A(n14246), .B(n13207), .C(n12666), .D(n14179), 
        .Z(n14278) );
  HS65_LL_NOR4ABX2 U13568 ( .A(n13202), .B(n13833), .C(n14164), .D(n14278), 
        .Z(n11389) );
  HS65_LL_NAND4ABX3 U13569 ( .A(n12668), .B(n14261), .C(n14175), .D(n11389), 
        .Z(n11392) );
  HS65_LL_NOR2X2 U13570 ( .A(n11391), .B(n11390), .Z(n14279) );
  HS65_LL_MX41X4 U13571 ( .D0(n11395), .S0(n14285), .D1(n11394), .S1(n14283), 
        .D2(n11393), .S2(n14281), .D3(n11392), .S3(n14279), .Z(n15432) );
  HS65_LL_IVX2 U13572 ( .A(sa10[1]), .Z(n13137) );
  HS65_LL_NOR2X2 U13573 ( .A(sa10[7]), .B(n13137), .Z(n14197) );
  HS65_LL_IVX2 U13574 ( .A(sa10[6]), .Z(n11985) );
  HS65_LL_NAND2X2 U13575 ( .A(n14197), .B(n11985), .Z(n11978) );
  HS65_LL_IVX2 U13576 ( .A(sa10[0]), .Z(n11396) );
  HS65_LL_NOR2X2 U13577 ( .A(sa10[3]), .B(n11396), .Z(n11407) );
  HS65_LL_NAND2X2 U13578 ( .A(sa10[5]), .B(n11407), .Z(n11401) );
  HS65_LL_NOR2X2 U13579 ( .A(n11978), .B(n11401), .Z(n13899) );
  HS65_LL_NAND3X2 U13580 ( .A(sa10[7]), .B(n11985), .C(n13137), .Z(n11418) );
  HS65_LL_NOR2X2 U13581 ( .A(n11418), .B(n11401), .Z(n14219) );
  HS65_LL_NAND2X2 U13582 ( .A(sa10[6]), .B(n13137), .Z(n11996) );
  HS65_LL_NAND3X2 U13583 ( .A(sa10[5]), .B(sa10[0]), .C(sa10[3]), .Z(n11979)
         );
  HS65_LL_NOR2X2 U13584 ( .A(n11996), .B(n11979), .Z(n11419) );
  HS65_LL_NAND2X2 U13585 ( .A(sa10[7]), .B(n11419), .Z(n13923) );
  HS65_LL_NAND2X2 U13586 ( .A(n11396), .B(sa10[3]), .Z(n11980) );
  HS65_LL_IVX2 U13587 ( .A(n11980), .Z(n11409) );
  HS65_LL_NAND2X2 U13588 ( .A(sa10[5]), .B(n11409), .Z(n13147) );
  HS65_LL_NAND2X2 U13589 ( .A(sa10[6]), .B(n14197), .Z(n11966) );
  HS65_LL_NOR2X2 U13590 ( .A(n13147), .B(n11966), .Z(n14211) );
  HS65_LL_NOR2AX3 U13591 ( .A(n13923), .B(n14211), .Z(n12111) );
  HS65_LL_NOR2X2 U13592 ( .A(sa10[7]), .B(n11996), .Z(n12103) );
  HS65_LL_NAND2X2 U13593 ( .A(n12103), .B(n11407), .Z(n12116) );
  HS65_LL_NOR2X2 U13594 ( .A(sa10[5]), .B(n12116), .Z(n12108) );
  HS65_LL_IVX2 U13595 ( .A(sa10[5]), .Z(n11964) );
  HS65_LL_NAND2X2 U13596 ( .A(n11409), .B(n11964), .Z(n12781) );
  HS65_LL_NOR2X2 U13597 ( .A(n12781), .B(n11966), .Z(n12102) );
  HS65_LL_IVX2 U13598 ( .A(n12102), .Z(n11968) );
  HS65_LL_NOR3X1 U13599 ( .A(sa10[6]), .B(sa10[7]), .C(sa10[1]), .Z(n11958) );
  HS65_LL_NOR2AX3 U13600 ( .A(n11958), .B(n11980), .Z(n13156) );
  HS65_LL_NAND2X2 U13601 ( .A(n13156), .B(n11964), .Z(n13916) );
  HS65_LL_NAND2X2 U13602 ( .A(n11968), .B(n13916), .Z(n12767) );
  HS65_LL_NAND3X2 U13603 ( .A(sa10[6]), .B(sa10[7]), .C(sa10[1]), .Z(n13146)
         );
  HS65_LL_IVX2 U13604 ( .A(n13146), .Z(n12120) );
  HS65_LL_NOR2X2 U13605 ( .A(sa10[0]), .B(sa10[3]), .Z(n11397) );
  HS65_LL_NAND2X2 U13606 ( .A(sa10[5]), .B(n11397), .Z(n11965) );
  HS65_LL_IVX2 U13607 ( .A(n11965), .Z(n14196) );
  HS65_LL_NAND2X2 U13608 ( .A(n12120), .B(n14196), .Z(n13924) );
  HS65_LL_NAND2X2 U13609 ( .A(n11407), .B(n11964), .Z(n11421) );
  HS65_LL_IVX2 U13610 ( .A(n11421), .Z(n11402) );
  HS65_LL_IVX2 U13611 ( .A(n11418), .Z(n11414) );
  HS65_LL_NAND2X2 U13612 ( .A(n11402), .B(n11414), .Z(n12772) );
  HS65_LL_NAND2X2 U13613 ( .A(n13924), .B(n12772), .Z(n14225) );
  HS65_LL_NOR3X1 U13614 ( .A(n12108), .B(n12767), .C(n14225), .Z(n11398) );
  HS65_LL_NAND4ABX3 U13615 ( .A(n13899), .B(n14219), .C(n12111), .D(n11398), 
        .Z(n13167) );
  HS65_LL_NOR3X1 U13616 ( .A(sa10[5]), .B(n11980), .C(n11418), .Z(n14889) );
  HS65_LL_NOR3X1 U13617 ( .A(sa10[5]), .B(sa10[0]), .C(sa10[3]), .Z(n11986) );
  HS65_LL_NAND3X2 U13618 ( .A(sa10[7]), .B(sa10[1]), .C(n11985), .Z(n11963) );
  HS65_LL_IVX2 U13619 ( .A(n11963), .Z(n12788) );
  HS65_LL_NAND2X2 U13620 ( .A(n11986), .B(n12788), .Z(n12761) );
  HS65_LL_IVX2 U13621 ( .A(n12761), .Z(n12127) );
  HS65_LL_NOR2X2 U13622 ( .A(n13147), .B(n11963), .Z(n13905) );
  HS65_LL_NOR3X1 U13623 ( .A(n14889), .B(n12127), .C(n13905), .Z(n11425) );
  HS65_LL_NAND2X2 U13624 ( .A(n11986), .B(n11414), .Z(n14190) );
  HS65_LL_IVX2 U13625 ( .A(n11978), .Z(n11406) );
  HS65_LL_NAND2X2 U13626 ( .A(n11406), .B(n11402), .Z(n14188) );
  HS65_LL_IVX2 U13627 ( .A(n13147), .Z(n13138) );
  HS65_LL_NAND3X2 U13628 ( .A(sa10[6]), .B(sa10[7]), .C(n13138), .Z(n12115) );
  HS65_LL_NOR2X2 U13629 ( .A(sa10[1]), .B(n12115), .Z(n13148) );
  HS65_LL_NAND2X2 U13630 ( .A(n11406), .B(n11986), .Z(n11960) );
  HS65_LL_IVX2 U13631 ( .A(n11960), .Z(n14872) );
  HS65_LL_NOR4ABX2 U13632 ( .A(n14190), .B(n14188), .C(n13148), .D(n14872), 
        .Z(n14883) );
  HS65_LL_NAND2X2 U13633 ( .A(n11425), .B(n14883), .Z(n14870) );
  HS65_LL_NOR2AX3 U13634 ( .A(n11419), .B(sa10[7]), .Z(n13164) );
  HS65_LL_IVX2 U13635 ( .A(n11401), .Z(n12119) );
  HS65_LL_NAND2X2 U13636 ( .A(n11958), .B(n12119), .Z(n12760) );
  HS65_LL_NAND2X2 U13637 ( .A(n11986), .B(n12120), .Z(n11995) );
  HS65_LL_NAND2X2 U13638 ( .A(n12760), .B(n11995), .Z(n11411) );
  HS65_LL_NOR2X2 U13639 ( .A(n13164), .B(n11411), .Z(n11959) );
  HS65_LL_AND2X4 U13640 ( .A(sa10[3]), .B(sa10[0]), .Z(n12132) );
  HS65_LL_NAND2X2 U13641 ( .A(n11964), .B(n12132), .Z(n11408) );
  HS65_LL_NAND3X2 U13642 ( .A(sa10[7]), .B(sa10[6]), .C(n13137), .Z(n11413) );
  HS65_LL_NOR2X2 U13643 ( .A(n11408), .B(n11413), .Z(n14209) );
  HS65_LL_AOI12X2 U13644 ( .A(n12119), .B(n12120), .C(n14209), .Z(n14223) );
  HS65_LL_NAND2X2 U13645 ( .A(n11958), .B(n14196), .Z(n12128) );
  HS65_LL_NOR3X1 U13646 ( .A(sa10[6]), .B(sa10[1]), .C(n11408), .Z(n14201) );
  HS65_LL_NOR2X2 U13647 ( .A(n11979), .B(n11418), .Z(n12777) );
  HS65_LL_NOR4ABX2 U13648 ( .A(n14223), .B(n12128), .C(n14201), .D(n12777), 
        .Z(n11399) );
  HS65_LL_NOR2X2 U13649 ( .A(n13146), .B(n11979), .Z(n13904) );
  HS65_LL_IVX2 U13650 ( .A(n11408), .Z(n11962) );
  HS65_LL_AND2X4 U13651 ( .A(n14197), .B(n11962), .Z(n12795) );
  HS65_LL_NOR2AX3 U13652 ( .A(n12795), .B(sa10[6]), .Z(n13903) );
  HS65_LL_NOR4ABX2 U13653 ( .A(n11959), .B(n11399), .C(n13904), .D(n13903), 
        .Z(n14203) );
  HS65_LL_NAND2X2 U13654 ( .A(sa10[6]), .B(sa10[7]), .Z(n11400) );
  HS65_LL_NOR2X2 U13655 ( .A(n11400), .B(n11421), .Z(n12751) );
  HS65_LL_NAND2X2 U13656 ( .A(sa10[1]), .B(n12751), .Z(n14861) );
  HS65_LL_NOR2X2 U13657 ( .A(n11965), .B(n11963), .Z(n12784) );
  HS65_LL_NOR2X2 U13658 ( .A(n11966), .B(n11401), .Z(n12758) );
  HS65_LL_IVX2 U13659 ( .A(n12758), .Z(n11984) );
  HS65_LL_NAND2X2 U13660 ( .A(n11402), .B(n12788), .Z(n12770) );
  HS65_LL_NAND2X2 U13661 ( .A(n11984), .B(n12770), .Z(n11403) );
  HS65_LL_NOR4ABX2 U13662 ( .A(n14203), .B(n14861), .C(n12784), .D(n11403), 
        .Z(n11426) );
  HS65_LL_OR2X4 U13663 ( .A(n12116), .B(n11964), .Z(n12756) );
  HS65_LL_NOR2X2 U13664 ( .A(n11421), .B(n11413), .Z(n12780) );
  HS65_LL_AOI12X2 U13665 ( .A(n12788), .B(n12119), .C(n12780), .Z(n11422) );
  HS65_LL_IVX2 U13666 ( .A(n11413), .Z(n11415) );
  HS65_LL_NAND2X2 U13667 ( .A(n11986), .B(n11415), .Z(n12789) );
  HS65_LL_IVX2 U13668 ( .A(n12789), .Z(n12134) );
  HS65_LL_NAND3X2 U13669 ( .A(n11985), .B(n14197), .C(n14196), .Z(n12131) );
  HS65_LL_IVX2 U13670 ( .A(n11979), .Z(n11405) );
  HS65_LL_NAND2X2 U13671 ( .A(n11406), .B(n11405), .Z(n12117) );
  HS65_LL_NAND2X2 U13672 ( .A(sa10[6]), .B(n12795), .Z(n13915) );
  HS65_LL_NAND3X2 U13673 ( .A(n12131), .B(n12117), .C(n13915), .Z(n14213) );
  HS65_LL_NOR4ABX2 U13674 ( .A(n12756), .B(n11422), .C(n12134), .D(n14213), 
        .Z(n11404) );
  HS65_LL_NAND4ABX3 U13675 ( .A(n13167), .B(n14870), .C(n11426), .D(n11404), 
        .Z(n11432) );
  HS65_LL_IVX2 U13676 ( .A(sa10[4]), .Z(n11428) );
  HS65_LL_NAND2X2 U13677 ( .A(sa10[2]), .B(n11428), .Z(n12774) );
  HS65_LL_IVX2 U13678 ( .A(n12774), .Z(n14899) );
  HS65_LL_NAND2X2 U13679 ( .A(n11962), .B(n12120), .Z(n13913) );
  HS65_LL_NAND2X2 U13680 ( .A(n13913), .B(n14190), .Z(n12765) );
  HS65_LL_NAND2X2 U13681 ( .A(sa10[7]), .B(n14201), .Z(n13162) );
  HS65_LL_NAND2X2 U13682 ( .A(n13162), .B(n14861), .Z(n12790) );
  HS65_LL_NOR2X2 U13683 ( .A(n13905), .B(n12790), .Z(n11972) );
  HS65_LL_NOR2X2 U13684 ( .A(n11978), .B(n12781), .Z(n12750) );
  HS65_LL_NOR2X2 U13685 ( .A(n11966), .B(n11979), .Z(n12114) );
  HS65_LL_NOR2X2 U13686 ( .A(n12781), .B(n11963), .Z(n12799) );
  HS65_LL_NOR3X1 U13687 ( .A(n12750), .B(n12114), .C(n12799), .Z(n13900) );
  HS65_LL_NAND3AX3 U13688 ( .A(n12765), .B(n11972), .C(n13900), .Z(n12786) );
  HS65_LL_NAND2X2 U13689 ( .A(n11958), .B(n11405), .Z(n12105) );
  HS65_LL_IVX2 U13690 ( .A(n12105), .Z(n12759) );
  HS65_LL_NAND2X2 U13691 ( .A(n12103), .B(n13138), .Z(n14886) );
  HS65_LL_NAND2X2 U13692 ( .A(n11406), .B(n13138), .Z(n13151) );
  HS65_LL_NAND4ABX3 U13693 ( .A(n12759), .B(n14872), .C(n14886), .D(n13151), 
        .Z(n14202) );
  HS65_LL_NAND2X2 U13694 ( .A(n14197), .B(n11986), .Z(n12764) );
  HS65_LL_NOR2X2 U13695 ( .A(n11985), .B(n12764), .Z(n11975) );
  HS65_LL_NOR2X2 U13696 ( .A(n13899), .B(n11975), .Z(n12110) );
  HS65_LL_NAND2X2 U13697 ( .A(n11968), .B(n12128), .Z(n12798) );
  HS65_LL_NAND2X2 U13698 ( .A(n11958), .B(n13138), .Z(n11989) );
  HS65_LL_NAND2X2 U13699 ( .A(n11989), .B(n12772), .Z(n14195) );
  HS65_LL_NAND2X2 U13700 ( .A(n11958), .B(n11407), .Z(n12769) );
  HS65_LL_NOR2X2 U13701 ( .A(sa10[5]), .B(n12769), .Z(n14864) );
  HS65_LL_NOR2X2 U13702 ( .A(n11408), .B(n11963), .Z(n12101) );
  HS65_LL_NOR2X2 U13703 ( .A(n14864), .B(n12101), .Z(n12122) );
  HS65_LL_NAND2X2 U13704 ( .A(n12756), .B(n12770), .Z(n13911) );
  HS65_LL_AOI112X2 U13705 ( .A(n12120), .B(n11409), .C(n14889), .D(n13911), 
        .Z(n11410) );
  HS65_LL_NAND4ABX3 U13706 ( .A(n12798), .B(n14195), .C(n12122), .D(n11410), 
        .Z(n13919) );
  HS65_LL_AOI112X2 U13707 ( .A(n12132), .B(n11415), .C(n11411), .D(n13919), 
        .Z(n11412) );
  HS65_LL_NAND4ABX3 U13708 ( .A(n12786), .B(n14202), .C(n12110), .D(n11412), 
        .Z(n11431) );
  HS65_LL_NOR2X2 U13709 ( .A(sa10[4]), .B(sa10[2]), .Z(n14891) );
  HS65_LL_NOR2AX3 U13710 ( .A(n14201), .B(sa10[7]), .Z(n14863) );
  HS65_LL_NAND4ABX3 U13711 ( .A(n13905), .B(n14863), .C(n13913), .D(n11995), 
        .Z(n13163) );
  HS65_LL_NAND2AX4 U13712 ( .A(n13163), .B(n13916), .Z(n13139) );
  HS65_LL_NAND2X2 U13713 ( .A(n11962), .B(n12103), .Z(n14198) );
  HS65_LL_IVX2 U13714 ( .A(n12784), .Z(n12794) );
  HS65_LL_NAND2X2 U13715 ( .A(n14198), .B(n12794), .Z(n12121) );
  HS65_LL_NOR2X2 U13716 ( .A(n12781), .B(n13146), .Z(n14210) );
  HS65_LL_IVX2 U13717 ( .A(n14210), .Z(n12104) );
  HS65_LL_NOR2X2 U13718 ( .A(n14219), .B(n14872), .Z(n12129) );
  HS65_LL_NOR2X2 U13719 ( .A(n12781), .B(n11413), .Z(n13906) );
  HS65_LL_NOR2X2 U13720 ( .A(n13906), .B(n12108), .Z(n12771) );
  HS65_LL_NOR2AX3 U13721 ( .A(n13162), .B(n13904), .Z(n12109) );
  HS65_LL_NOR2X2 U13722 ( .A(n11965), .B(n11413), .Z(n11992) );
  HS65_LL_NAND2X2 U13723 ( .A(n14196), .B(n11414), .Z(n13912) );
  HS65_LL_NAND2X2 U13724 ( .A(n12119), .B(n11415), .Z(n14220) );
  HS65_LL_NAND3X2 U13725 ( .A(n12756), .B(n13912), .C(n14220), .Z(n11998) );
  HS65_LL_NOR3X1 U13726 ( .A(n12759), .B(n11992), .C(n11998), .Z(n11416) );
  HS65_LL_NAND3X2 U13727 ( .A(n12771), .B(n12109), .C(n11416), .Z(n14901) );
  HS65_LL_NOR4ABX2 U13728 ( .A(n11984), .B(n12760), .C(n14901), .D(n14213), 
        .Z(n11417) );
  HS65_LL_OAI21X2 U13729 ( .A(n11980), .B(n11418), .C(n11417), .Z(n13155) );
  HS65_LL_NOR4ABX2 U13730 ( .A(n12104), .B(n12129), .C(n13155), .D(n11419), 
        .Z(n11420) );
  HS65_LL_NAND4ABX3 U13731 ( .A(n13139), .B(n12121), .C(n11420), .D(n14861), 
        .Z(n11430) );
  HS65_LL_NAND2X2 U13732 ( .A(sa10[4]), .B(sa10[2]), .Z(n14895) );
  HS65_LL_IVX2 U13733 ( .A(n14895), .Z(n14233) );
  HS65_LL_NOR2X2 U13734 ( .A(n12101), .B(n11992), .Z(n14215) );
  HS65_LL_NOR2X2 U13735 ( .A(n11966), .B(n11421), .Z(n14221) );
  HS65_LL_AOI12X2 U13736 ( .A(n12120), .B(n13138), .C(n14221), .Z(n11961) );
  HS65_LL_IVX2 U13737 ( .A(n14886), .Z(n12112) );
  HS65_LL_NOR4ABX2 U13738 ( .A(n11961), .B(n11422), .C(n12112), .D(n12767), 
        .Z(n11424) );
  HS65_LL_NOR2X2 U13739 ( .A(sa10[6]), .B(sa10[1]), .Z(n11423) );
  HS65_LL_NAND3X2 U13740 ( .A(sa10[7]), .B(n11423), .C(n13138), .Z(n14212) );
  HS65_LL_NAND3X2 U13741 ( .A(n11424), .B(n14212), .C(n14188), .Z(n13921) );
  HS65_LL_NAND3X2 U13742 ( .A(n11425), .B(n12104), .C(n13912), .Z(n14884) );
  HS65_LL_NOR3AX2 U13743 ( .A(n11426), .B(n13921), .C(n14884), .Z(n11427) );
  HS65_LL_NAND3X2 U13744 ( .A(n14215), .B(n11427), .C(n11989), .Z(n11429) );
  HS65_LL_NOR2X2 U13745 ( .A(sa10[2]), .B(n11428), .Z(n14893) );
  HS65_LL_MX41X4 U13746 ( .D0(n11432), .S0(n14899), .D1(n11431), .S1(n14891), 
        .D2(n11430), .S2(n14233), .D3(n11429), .S3(n14893), .Z(n15342) );
  HS65_LL_IVX2 U13747 ( .A(sa32[6]), .Z(n13278) );
  HS65_LL_IVX2 U13748 ( .A(sa32[7]), .Z(n13277) );
  HS65_LL_NAND3X2 U13749 ( .A(sa32[1]), .B(n13278), .C(n13277), .Z(n13189) );
  HS65_LL_NAND2X2 U13750 ( .A(sa32[3]), .B(sa32[0]), .Z(n11496) );
  HS65_LL_NOR2X2 U13751 ( .A(sa32[5]), .B(n11496), .Z(n11475) );
  HS65_LL_IVX2 U13752 ( .A(n11475), .Z(n11456) );
  HS65_LL_NOR2X2 U13753 ( .A(n13189), .B(n11456), .Z(n13180) );
  HS65_LL_IVX2 U13754 ( .A(sa32[0]), .Z(n11437) );
  HS65_LL_NOR2X2 U13755 ( .A(sa32[3]), .B(n11437), .Z(n12087) );
  HS65_LL_IVX2 U13756 ( .A(sa32[5]), .Z(n11434) );
  HS65_LL_NAND2X2 U13757 ( .A(n12087), .B(n11434), .Z(n11459) );
  HS65_LL_IVX2 U13758 ( .A(n11459), .Z(n11446) );
  HS65_LL_NOR3X1 U13759 ( .A(sa32[6]), .B(sa32[1]), .C(n13277), .Z(n11438) );
  HS65_LL_NAND2X2 U13760 ( .A(n11446), .B(n11438), .Z(n11468) );
  HS65_LL_NAND2X2 U13761 ( .A(sa32[1]), .B(n13277), .Z(n11457) );
  HS65_LL_NOR2X2 U13762 ( .A(n13278), .B(n11457), .Z(n11447) );
  HS65_LL_NOR3X1 U13763 ( .A(sa32[3]), .B(sa32[0]), .C(n11434), .Z(n13271) );
  HS65_LL_NAND2X2 U13764 ( .A(n11447), .B(n13271), .Z(n13193) );
  HS65_LL_NAND2X2 U13765 ( .A(n11468), .B(n13193), .Z(n14706) );
  HS65_LL_NAND2X2 U13766 ( .A(sa32[7]), .B(sa32[1]), .Z(n14723) );
  HS65_LL_IVX2 U13767 ( .A(n14723), .Z(n13270) );
  HS65_LL_NAND2X2 U13768 ( .A(n13270), .B(n13278), .Z(n11444) );
  HS65_LL_IVX2 U13769 ( .A(n11444), .Z(n13727) );
  HS65_LL_NAND2X2 U13770 ( .A(n13727), .B(n11475), .Z(n11472) );
  HS65_LL_IVX2 U13771 ( .A(n11472), .Z(n13247) );
  HS65_LL_NOR3X2 U13772 ( .A(sa32[6]), .B(sa32[7]), .C(sa32[1]), .Z(n12086) );
  HS65_LL_NAND2X2 U13773 ( .A(n12086), .B(n13271), .Z(n11497) );
  HS65_LL_NAND2X2 U13774 ( .A(sa32[5]), .B(n12087), .Z(n11492) );
  HS65_LL_IVX2 U13775 ( .A(n11492), .Z(n11450) );
  HS65_LL_NAND2X2 U13776 ( .A(n11438), .B(n11450), .Z(n11487) );
  HS65_LL_NAND2X2 U13777 ( .A(n11497), .B(n11487), .Z(n14346) );
  HS65_LL_NOR2X2 U13778 ( .A(n13247), .B(n14346), .Z(n12088) );
  HS65_LL_NOR2AX3 U13779 ( .A(sa32[3]), .B(sa32[0]), .Z(n14733) );
  HS65_LL_NAND2X2 U13780 ( .A(n14733), .B(n11434), .Z(n14722) );
  HS65_LL_IVX2 U13781 ( .A(n14722), .Z(n13729) );
  HS65_LL_AND2X4 U13782 ( .A(n11447), .B(n13729), .Z(n11491) );
  HS65_LL_NAND2X2 U13783 ( .A(n12086), .B(n11450), .Z(n11476) );
  HS65_LL_NOR3X1 U13784 ( .A(sa32[5]), .B(sa32[3]), .C(sa32[0]), .Z(n12056) );
  HS65_LL_NOR3X1 U13785 ( .A(n13278), .B(sa32[7]), .C(sa32[1]), .Z(n11477) );
  HS65_LL_NAND2X2 U13786 ( .A(n12056), .B(n11477), .Z(n14728) );
  HS65_LL_NAND2X2 U13787 ( .A(n11476), .B(n14728), .Z(n13289) );
  HS65_LL_NAND2X2 U13788 ( .A(n11446), .B(n12086), .Z(n13248) );
  HS65_LL_NAND2X2 U13789 ( .A(n13729), .B(n12086), .Z(n14348) );
  HS65_LL_NAND2X2 U13790 ( .A(n13248), .B(n14348), .Z(n12064) );
  HS65_LL_NAND2X2 U13791 ( .A(n11438), .B(n12056), .Z(n14729) );
  HS65_LL_IVX2 U13792 ( .A(n12056), .Z(n13282) );
  HS65_LL_NOR2X2 U13793 ( .A(n13189), .B(n13282), .Z(n14735) );
  HS65_LL_NOR2AX3 U13794 ( .A(n14729), .B(n14735), .Z(n11489) );
  HS65_LL_NAND2X2 U13795 ( .A(sa32[6]), .B(n13270), .Z(n11493) );
  HS65_LL_IVX2 U13796 ( .A(n11493), .Z(n11442) );
  HS65_LL_NAND2X2 U13797 ( .A(n11442), .B(n13271), .Z(n13739) );
  HS65_LL_NAND4ABX3 U13798 ( .A(n13289), .B(n12064), .C(n11489), .D(n13739), 
        .Z(n11433) );
  HS65_LL_NOR2X2 U13799 ( .A(n11493), .B(n11456), .Z(n13741) );
  HS65_LL_NAND2X2 U13800 ( .A(sa32[5]), .B(n14733), .Z(n13188) );
  HS65_LL_NOR3X1 U13801 ( .A(sa32[1]), .B(n13277), .C(n13278), .Z(n11474) );
  HS65_LL_IVX2 U13802 ( .A(n11474), .Z(n11458) );
  HS65_LL_NOR2X2 U13803 ( .A(n13188), .B(n11458), .Z(n13752) );
  HS65_LL_NOR2X2 U13804 ( .A(n13741), .B(n13752), .Z(n11460) );
  HS65_LL_NAND2X2 U13805 ( .A(n11447), .B(n12056), .Z(n14357) );
  HS65_LL_NAND4ABX3 U13806 ( .A(n11491), .B(n11433), .C(n11460), .D(n14357), 
        .Z(n13750) );
  HS65_LL_NOR2X2 U13807 ( .A(n11434), .B(n11496), .Z(n13728) );
  HS65_LL_IVX2 U13808 ( .A(n13728), .Z(n12055) );
  HS65_LL_NOR2X2 U13809 ( .A(n12055), .B(n11493), .Z(n13257) );
  HS65_LL_NOR2X2 U13810 ( .A(n14722), .B(n13189), .Z(n12084) );
  HS65_LL_IVX2 U13811 ( .A(n12084), .Z(n13279) );
  HS65_LL_NOR2X2 U13812 ( .A(n14722), .B(n11493), .Z(n11503) );
  HS65_LL_IVX2 U13813 ( .A(n11503), .Z(n13254) );
  HS65_LL_IVX2 U13814 ( .A(n13188), .Z(n11478) );
  HS65_LL_NAND2X2 U13815 ( .A(n11447), .B(n11478), .Z(n14364) );
  HS65_LL_NAND3X2 U13816 ( .A(n13279), .B(n13254), .C(n14364), .Z(n13735) );
  HS65_LL_NOR2X2 U13817 ( .A(n11493), .B(n11459), .Z(n11485) );
  HS65_LL_IVX2 U13818 ( .A(n12086), .Z(n11435) );
  HS65_LL_NAND2X2 U13819 ( .A(n11475), .B(n11477), .Z(n13178) );
  HS65_LL_OAI21X2 U13820 ( .A(n11435), .B(n13282), .C(n13178), .Z(n14731) );
  HS65_LL_NOR2X2 U13821 ( .A(n11485), .B(n14731), .Z(n11454) );
  HS65_LL_IVX2 U13822 ( .A(n13189), .Z(n14732) );
  HS65_LL_NAND2X2 U13823 ( .A(n14732), .B(n13271), .Z(n14360) );
  HS65_LL_AND2X4 U13824 ( .A(n11454), .B(n14360), .Z(n13252) );
  HS65_LL_NOR2X2 U13825 ( .A(n11459), .B(n11458), .Z(n12071) );
  HS65_LL_IVX2 U13826 ( .A(n12071), .Z(n14366) );
  HS65_LL_NAND4ABX3 U13827 ( .A(n13257), .B(n13735), .C(n13252), .D(n14366), 
        .Z(n13177) );
  HS65_LL_NOR2X2 U13828 ( .A(n11456), .B(n11435), .Z(n14700) );
  HS65_LL_NAND2X2 U13829 ( .A(n13727), .B(n11446), .Z(n14372) );
  HS65_LL_NOR3X1 U13830 ( .A(sa32[1]), .B(n13278), .C(n14722), .Z(n13256) );
  HS65_LL_NAND2X2 U13831 ( .A(sa32[7]), .B(n13256), .Z(n12076) );
  HS65_LL_NAND2X2 U13832 ( .A(n14372), .B(n12076), .Z(n13758) );
  HS65_LL_NAND2X2 U13833 ( .A(n11446), .B(n11477), .Z(n11490) );
  HS65_LL_NAND2X2 U13834 ( .A(n11477), .B(n13271), .Z(n14709) );
  HS65_LL_NAND4ABX3 U13835 ( .A(n14700), .B(n13758), .C(n11490), .D(n14709), 
        .Z(n13292) );
  HS65_LL_NOR3X1 U13836 ( .A(n13750), .B(n13177), .C(n13292), .Z(n11436) );
  HS65_LL_NAND4ABX3 U13837 ( .A(n13180), .B(n14706), .C(n12088), .D(n11436), 
        .Z(n11466) );
  HS65_LL_IVX2 U13838 ( .A(sa32[2]), .Z(n11441) );
  HS65_LL_NOR2X2 U13839 ( .A(sa32[4]), .B(n11441), .Z(n14748) );
  HS65_LL_NAND3X2 U13840 ( .A(sa32[5]), .B(sa32[3]), .C(n14732), .Z(n12082) );
  HS65_LL_NOR2X2 U13841 ( .A(n11437), .B(n12082), .Z(n14355) );
  HS65_LL_IVX2 U13842 ( .A(n11438), .Z(n12054) );
  HS65_LL_NOR2X2 U13843 ( .A(n14722), .B(n12054), .Z(n13263) );
  HS65_LL_NAND2X2 U13844 ( .A(n11478), .B(n12086), .Z(n14703) );
  HS65_LL_NAND2AX4 U13845 ( .A(n13263), .B(n14703), .Z(n11470) );
  HS65_LL_NAND2X2 U13846 ( .A(n11475), .B(n11438), .Z(n14701) );
  HS65_LL_IVX2 U13847 ( .A(n14701), .Z(n13181) );
  HS65_LL_AOI12X2 U13848 ( .A(n13256), .B(n13277), .C(n13181), .Z(n11452) );
  HS65_LL_AOI12X2 U13849 ( .A(n11438), .B(n13728), .C(n11491), .Z(n13255) );
  HS65_LL_NAND4ABX3 U13850 ( .A(n14355), .B(n11470), .C(n11452), .D(n13255), 
        .Z(n13284) );
  HS65_LL_NAND2X2 U13851 ( .A(n13728), .B(n12086), .Z(n14736) );
  HS65_LL_NAND2X2 U13852 ( .A(n11477), .B(n11450), .Z(n11481) );
  HS65_LL_IVX2 U13853 ( .A(n11481), .Z(n13759) );
  HS65_LL_NAND2X2 U13854 ( .A(n13728), .B(n11477), .Z(n12067) );
  HS65_LL_IVX2 U13855 ( .A(n12067), .Z(n11494) );
  HS65_LL_AND2X4 U13856 ( .A(n13271), .B(n11438), .Z(n11502) );
  HS65_LL_NOR2X2 U13857 ( .A(n11494), .B(n11502), .Z(n13719) );
  HS65_LL_NAND2X2 U13858 ( .A(n11447), .B(n11450), .Z(n12051) );
  HS65_LL_NAND3X2 U13859 ( .A(n13719), .B(n13248), .C(n12051), .Z(n11439) );
  HS65_LL_NOR3AX2 U13860 ( .A(n14736), .B(n13759), .C(n11439), .Z(n14724) );
  HS65_LL_NOR2X2 U13861 ( .A(n12055), .B(n11444), .Z(n12080) );
  HS65_LL_NAND3X2 U13862 ( .A(n13278), .B(n13270), .C(n13271), .Z(n13717) );
  HS65_LL_IVX2 U13863 ( .A(n13717), .Z(n12075) );
  HS65_LL_NOR3X1 U13864 ( .A(n12080), .B(n13180), .C(n12075), .Z(n12070) );
  HS65_LL_NAND2X2 U13865 ( .A(n14732), .B(n11450), .Z(n13731) );
  HS65_LL_NOR2X2 U13866 ( .A(n11444), .B(n13282), .Z(n13737) );
  HS65_LL_NOR4ABX2 U13867 ( .A(n12070), .B(n13731), .C(n13737), .D(n13289), 
        .Z(n11440) );
  HS65_LL_NAND4ABX3 U13868 ( .A(n13177), .B(n13284), .C(n14724), .D(n11440), 
        .Z(n11465) );
  HS65_LL_NAND2X2 U13869 ( .A(sa32[4]), .B(n11441), .Z(n13744) );
  HS65_LL_IVX2 U13870 ( .A(n13744), .Z(n14746) );
  HS65_LL_NOR4ABX2 U13871 ( .A(n13717), .B(n14709), .C(n13257), .D(n13256), 
        .Z(n11449) );
  HS65_LL_IVX2 U13872 ( .A(n11476), .Z(n13753) );
  HS65_LL_NOR2X2 U13873 ( .A(n13263), .B(n13753), .Z(n11483) );
  HS65_LL_AOI12X2 U13874 ( .A(n12086), .B(n12056), .C(n11494), .Z(n13264) );
  HS65_LL_NAND2X2 U13875 ( .A(n11442), .B(n12056), .Z(n12077) );
  HS65_LL_OAI21X2 U13876 ( .A(n13188), .B(n13189), .C(n12077), .Z(n11479) );
  HS65_LL_NAND2X2 U13877 ( .A(n13271), .B(n11474), .Z(n13722) );
  HS65_LL_NAND2X2 U13878 ( .A(n11472), .B(n13722), .Z(n14740) );
  HS65_LL_NOR4ABX2 U13879 ( .A(n11483), .B(n13264), .C(n11479), .D(n14740), 
        .Z(n13186) );
  HS65_LL_NAND2X2 U13880 ( .A(n11468), .B(n13739), .Z(n14712) );
  HS65_LL_OAI21X2 U13881 ( .A(n12054), .B(n12055), .C(n13731), .Z(n11451) );
  HS65_LL_NOR2X2 U13882 ( .A(n11492), .B(n11458), .Z(n13269) );
  HS65_LL_NAND2X2 U13883 ( .A(n11447), .B(n11475), .Z(n13716) );
  HS65_LL_NAND3AX3 U13884 ( .A(n13269), .B(n14736), .C(n13716), .Z(n11443) );
  HS65_LL_NOR3X1 U13885 ( .A(n14712), .B(n11451), .C(n11443), .Z(n13175) );
  HS65_LL_NOR2X2 U13886 ( .A(n11444), .B(n13188), .Z(n12062) );
  HS65_LL_NOR2X2 U13887 ( .A(n12062), .B(n11485), .Z(n13757) );
  HS65_LL_NAND2X2 U13888 ( .A(n13728), .B(n11447), .Z(n13266) );
  HS65_LL_NAND2X2 U13889 ( .A(n13757), .B(n13266), .Z(n12089) );
  HS65_LL_NAND2X2 U13890 ( .A(n13729), .B(n13727), .Z(n13718) );
  HS65_LL_NAND2AX4 U13891 ( .A(n13741), .B(n13718), .Z(n13751) );
  HS65_LL_NOR3X1 U13892 ( .A(n12084), .B(n12089), .C(n13751), .Z(n11445) );
  HS65_LL_NAND3X2 U13893 ( .A(n11445), .B(n14701), .C(n14729), .Z(n12068) );
  HS65_LL_NOR2X2 U13894 ( .A(n13188), .B(n11493), .Z(n11504) );
  HS65_LL_NAND2X2 U13895 ( .A(n11447), .B(n11446), .Z(n13179) );
  HS65_LL_IVX2 U13896 ( .A(n13179), .Z(n14708) );
  HS65_LL_NOR2X2 U13897 ( .A(n12071), .B(n14708), .Z(n11505) );
  HS65_LL_NAND4ABX3 U13898 ( .A(n11504), .B(n14735), .C(n11505), .D(n14703), 
        .Z(n14727) );
  HS65_LL_NOR4ABX2 U13899 ( .A(n13186), .B(n13175), .C(n12068), .D(n14727), 
        .Z(n11448) );
  HS65_LL_NAND3X2 U13900 ( .A(n11449), .B(n11448), .C(n14364), .Z(n11464) );
  HS65_LL_NAND2X2 U13901 ( .A(sa32[4]), .B(sa32[2]), .Z(n14380) );
  HS65_LL_IVX2 U13902 ( .A(n14380), .Z(n14744) );
  HS65_LL_NAND2X2 U13903 ( .A(n12056), .B(n11474), .Z(n14361) );
  HS65_LL_NAND2X2 U13904 ( .A(n14361), .B(n13193), .Z(n12073) );
  HS65_LL_NAND2X2 U13905 ( .A(n13727), .B(n11450), .Z(n14710) );
  HS65_LL_NOR4ABX2 U13906 ( .A(n11452), .B(n14710), .C(n12080), .D(n11451), 
        .Z(n11453) );
  HS65_LL_NAND4ABX3 U13907 ( .A(n14708), .B(n12073), .C(n11454), .D(n11453), 
        .Z(n13725) );
  HS65_LL_NAND2X2 U13908 ( .A(n13279), .B(n11497), .Z(n12063) );
  HS65_LL_NOR2X2 U13909 ( .A(sa32[1]), .B(n13277), .Z(n11455) );
  HS65_LL_NAND2X2 U13910 ( .A(n11478), .B(n11455), .Z(n13173) );
  HS65_LL_NOR2X2 U13911 ( .A(sa32[6]), .B(n13173), .Z(n13287) );
  HS65_LL_NOR2X2 U13912 ( .A(n11491), .B(n13287), .Z(n11506) );
  HS65_LL_NOR2X2 U13913 ( .A(n11457), .B(n11456), .Z(n13275) );
  HS65_LL_NAND2X2 U13914 ( .A(n11487), .B(n14364), .Z(n13286) );
  HS65_LL_NOR2X2 U13915 ( .A(n13275), .B(n13286), .Z(n13743) );
  HS65_LL_NOR2X2 U13916 ( .A(n12055), .B(n11458), .Z(n13740) );
  HS65_LL_NOR2X2 U13917 ( .A(n14735), .B(n13740), .Z(n11488) );
  HS65_LL_IVX2 U13918 ( .A(n11490), .Z(n12050) );
  HS65_LL_NOR2X2 U13919 ( .A(n13759), .B(n11504), .Z(n11469) );
  HS65_LL_NOR2X2 U13920 ( .A(n13189), .B(n11459), .Z(n13258) );
  HS65_LL_IVX2 U13921 ( .A(n12051), .Z(n11499) );
  HS65_LL_NOR3AX2 U13922 ( .A(n13266), .B(n13258), .C(n11499), .Z(n13274) );
  HS65_LL_NAND3X2 U13923 ( .A(n11469), .B(n11460), .C(n13274), .Z(n11461) );
  HS65_LL_NOR3X1 U13924 ( .A(n13737), .B(n12050), .C(n11461), .Z(n14352) );
  HS65_LL_NAND3X2 U13925 ( .A(n11488), .B(n14352), .C(n14360), .Z(n14716) );
  HS65_LL_NOR4ABX2 U13926 ( .A(n13743), .B(n13718), .C(n12075), .D(n14716), 
        .Z(n11462) );
  HS65_LL_NAND4ABX3 U13927 ( .A(n13725), .B(n12063), .C(n11506), .D(n11462), 
        .Z(n11463) );
  HS65_LL_NOR2X2 U13928 ( .A(sa32[4]), .B(sa32[2]), .Z(n14742) );
  HS65_LL_MX41X4 U13929 ( .D0(n11466), .S0(n14748), .D1(n11465), .S1(n14746), 
        .D2(n11464), .S2(n14744), .D3(n11463), .S3(n14742), .Z(n15519) );
  HS65_LL_MUXI21X2 U13930 ( .D0(n11559), .D1(w3[10]), .S0(n15519), .Z(n11467)
         );
  HS65_LLS_XOR3X2 U13931 ( .A(n15432), .B(n15342), .C(n11467), .Z(n11562) );
  HS65_LL_NAND2X2 U13932 ( .A(n14372), .B(n11497), .Z(n13191) );
  HS65_LL_NAND4ABX3 U13933 ( .A(n11470), .B(n13191), .C(n11469), .D(n11468), 
        .Z(n11471) );
  HS65_LL_NOR3X1 U13934 ( .A(n11491), .B(n11503), .C(n11471), .Z(n11473) );
  HS65_LL_NAND3X2 U13935 ( .A(n11473), .B(n13248), .C(n11472), .Z(n13726) );
  HS65_LL_NAND2X2 U13936 ( .A(n11475), .B(n11474), .Z(n14720) );
  HS65_LL_NAND2X2 U13937 ( .A(n14720), .B(n11476), .Z(n14711) );
  HS65_LL_NAND2X2 U13938 ( .A(n11478), .B(n11477), .Z(n14371) );
  HS65_LL_NAND2X2 U13939 ( .A(n14736), .B(n14357), .Z(n12091) );
  HS65_LL_NOR4ABX2 U13940 ( .A(n14371), .B(n13731), .C(n12091), .D(n11479), 
        .Z(n11480) );
  HS65_LL_NAND4ABX3 U13941 ( .A(n13726), .B(n14711), .C(n11488), .D(n11480), 
        .Z(n11517) );
  HS65_LL_NAND2X2 U13942 ( .A(n14360), .B(n13716), .Z(n14719) );
  HS65_LL_NOR2X2 U13943 ( .A(n14355), .B(n14719), .Z(n14737) );
  HS65_LL_NAND2X2 U13944 ( .A(n14736), .B(n11490), .Z(n14368) );
  HS65_LL_NOR2X2 U13945 ( .A(n11502), .B(n13269), .Z(n14713) );
  HS65_LL_NAND2X2 U13946 ( .A(n14713), .B(n11481), .Z(n12083) );
  HS65_LL_NOR2X2 U13947 ( .A(n13181), .B(n13257), .Z(n14353) );
  HS65_LL_NAND3X2 U13948 ( .A(n14353), .B(n13722), .C(n12076), .Z(n11482) );
  HS65_LL_NOR3X1 U13949 ( .A(n14368), .B(n12083), .C(n11482), .Z(n13734) );
  HS65_LL_NAND3X2 U13950 ( .A(n14737), .B(n13734), .C(n11483), .Z(n11484) );
  HS65_LL_NOR3X1 U13951 ( .A(n11499), .B(n13287), .C(n11484), .Z(n13190) );
  HS65_LL_NAND2X2 U13952 ( .A(n13254), .B(n13178), .Z(n12079) );
  HS65_LL_IVX2 U13953 ( .A(n12077), .Z(n13276) );
  HS65_LL_NOR2X2 U13954 ( .A(n13276), .B(n14700), .Z(n11495) );
  HS65_LL_NOR2X2 U13955 ( .A(n12062), .B(n13741), .Z(n13721) );
  HS65_LL_NAND2X2 U13956 ( .A(n11495), .B(n13721), .Z(n14376) );
  HS65_LL_NOR2X2 U13957 ( .A(n11485), .B(n12075), .Z(n11500) );
  HS65_LL_NAND4ABX3 U13958 ( .A(n12079), .B(n14376), .C(n11500), .D(n14348), 
        .Z(n11486) );
  HS65_LL_NOR4ABX2 U13959 ( .A(n11488), .B(n11487), .C(n11486), .D(n11494), 
        .Z(n11515) );
  HS65_LL_NOR3X1 U13960 ( .A(n12062), .B(n13263), .C(n13737), .Z(n11508) );
  HS65_LL_NOR2X2 U13961 ( .A(n13258), .B(n13752), .Z(n12053) );
  HS65_LL_NAND3X2 U13962 ( .A(n11508), .B(n12053), .C(n11489), .Z(n13290) );
  HS65_LL_NAND4ABX3 U13963 ( .A(n13759), .B(n12071), .C(n14737), .D(n14710), 
        .Z(n11501) );
  HS65_LL_NAND2AX4 U13964 ( .A(n11491), .B(n11490), .Z(n12065) );
  HS65_LL_IVX2 U13965 ( .A(n13731), .Z(n12074) );
  HS65_LL_NOR3X1 U13966 ( .A(n13740), .B(n12074), .C(n13286), .Z(n14354) );
  HS65_LL_NAND4ABX3 U13967 ( .A(n12065), .B(n14712), .C(n14354), .D(n14348), 
        .Z(n13183) );
  HS65_LL_NOR2X2 U13968 ( .A(n11493), .B(n11492), .Z(n14707) );
  HS65_LL_NOR2AX3 U13969 ( .A(n11495), .B(n11494), .Z(n12061) );
  HS65_LL_NOR2X2 U13970 ( .A(n13257), .B(n13180), .Z(n13756) );
  HS65_LL_OA112X4 U13971 ( .A(n11496), .B(n12054), .C(n12061), .D(n13756), .Z(
        n11498) );
  HS65_LL_NAND4ABX3 U13972 ( .A(n14707), .B(n14711), .C(n11498), .D(n11497), 
        .Z(n14741) );
  HS65_LL_NOR4ABX2 U13973 ( .A(n11500), .B(n14372), .C(n11499), .D(n14741), 
        .Z(n11510) );
  HS65_LL_NAND4ABX3 U13974 ( .A(n11501), .B(n13183), .C(n11510), .D(n14361), 
        .Z(n11513) );
  HS65_LL_NOR2X2 U13975 ( .A(n11503), .B(n11502), .Z(n13288) );
  HS65_LL_NAND2X2 U13976 ( .A(n14371), .B(n14348), .Z(n14363) );
  HS65_LL_NAND2AX4 U13977 ( .A(n11504), .B(n14710), .Z(n13730) );
  HS65_LL_IVX2 U13978 ( .A(n13258), .Z(n14367) );
  HS65_LL_NAND3X2 U13979 ( .A(n11506), .B(n11505), .C(n14367), .Z(n11507) );
  HS65_LL_NOR3X1 U13980 ( .A(n14363), .B(n13730), .C(n11507), .Z(n13746) );
  HS65_LL_IVX2 U13981 ( .A(n11508), .Z(n11509) );
  HS65_LL_NOR4ABX2 U13982 ( .A(n11510), .B(n13746), .C(n11509), .D(n14740), 
        .Z(n11511) );
  HS65_LL_AOI13X2 U13983 ( .A(n13288), .B(n11511), .C(n14703), .D(n13744), .Z(
        n11512) );
  HS65_LL_CBI4I6X2 U13984 ( .A(n13290), .B(n11513), .C(n14748), .D(n11512), 
        .Z(n11514) );
  HS65_LL_CBI4I1X3 U13985 ( .A(n13190), .B(n11515), .C(n14380), .D(n11514), 
        .Z(n11516) );
  HS65_LL_CBI4I6X2 U13986 ( .A(n12068), .B(n11517), .C(n14742), .D(n11516), 
        .Z(n15518) );
  HS65_LL_IVX2 U13987 ( .A(sa03[1]), .Z(n11526) );
  HS65_LL_NOR2X2 U13988 ( .A(sa03[7]), .B(n11526), .Z(n11522) );
  HS65_LL_NAND2X2 U13989 ( .A(sa03[6]), .B(n11522), .Z(n12026) );
  HS65_LL_IVX2 U13990 ( .A(sa03[0]), .Z(n11521) );
  HS65_LL_NOR2X2 U13991 ( .A(sa03[3]), .B(n11521), .Z(n13114) );
  HS65_LL_NAND2X2 U13992 ( .A(sa03[5]), .B(n13114), .Z(n11540) );
  HS65_LL_NOR2X2 U13993 ( .A(n12026), .B(n11540), .Z(n15215) );
  HS65_LL_IVX2 U13994 ( .A(sa03[5]), .Z(n11528) );
  HS65_LL_NAND2X2 U13995 ( .A(n13114), .B(n11528), .Z(n12007) );
  HS65_LL_IVX2 U13996 ( .A(sa03[7]), .Z(n11518) );
  HS65_LL_NOR2X2 U13997 ( .A(sa03[6]), .B(n11518), .Z(n12695) );
  HS65_LL_NAND2X2 U13998 ( .A(sa03[1]), .B(n12695), .Z(n14594) );
  HS65_LL_NOR2X2 U13999 ( .A(n12007), .B(n14594), .Z(n13099) );
  HS65_LL_NAND2X2 U14000 ( .A(sa03[6]), .B(sa03[7]), .Z(n14574) );
  HS65_LL_NOR2X2 U14001 ( .A(sa03[1]), .B(n14574), .Z(n11548) );
  HS65_LL_NAND2X2 U14002 ( .A(sa03[0]), .B(sa03[3]), .Z(n12022) );
  HS65_LL_NOR2X2 U14003 ( .A(sa03[5]), .B(n12022), .Z(n13104) );
  HS65_LL_NAND2X2 U14004 ( .A(n11548), .B(n13104), .Z(n14592) );
  HS65_LL_NAND3X2 U14005 ( .A(sa03[1]), .B(sa03[6]), .C(sa03[7]), .Z(n11544)
         );
  HS65_LL_IVX2 U14006 ( .A(n11544), .Z(n11525) );
  HS65_LL_IVX2 U14007 ( .A(n11540), .Z(n11533) );
  HS65_LL_NAND2X2 U14008 ( .A(n11525), .B(n11533), .Z(n13773) );
  HS65_LL_NAND2X2 U14009 ( .A(n14592), .B(n13773), .Z(n14589) );
  HS65_LL_NAND2X2 U14010 ( .A(n11526), .B(n12695), .Z(n12027) );
  HS65_LL_IVX2 U14011 ( .A(n12027), .Z(n13105) );
  HS65_LL_NAND2X2 U14012 ( .A(n13105), .B(n13104), .Z(n12720) );
  HS65_LL_NOR2X2 U14013 ( .A(n11528), .B(n12022), .Z(n12714) );
  HS65_LL_NAND2X2 U14014 ( .A(n11525), .B(n12714), .Z(n14601) );
  HS65_LL_NAND2X2 U14015 ( .A(n12720), .B(n14601), .Z(n13774) );
  HS65_LL_IVX2 U14016 ( .A(sa03[6]), .Z(n12006) );
  HS65_LL_NAND3X2 U14017 ( .A(n11526), .B(n12006), .C(n11518), .Z(n13119) );
  HS65_LL_IVX2 U14018 ( .A(n13119), .Z(n13115) );
  HS65_LL_NAND2X2 U14019 ( .A(n13115), .B(n13104), .Z(n14607) );
  HS65_LL_NAND2X2 U14020 ( .A(n12714), .B(n13105), .Z(n13096) );
  HS65_LL_NAND2X2 U14021 ( .A(n14607), .B(n13096), .Z(n15222) );
  HS65_LL_NOR3X1 U14022 ( .A(n14589), .B(n13774), .C(n15222), .Z(n11519) );
  HS65_LL_NOR3X1 U14023 ( .A(sa03[0]), .B(sa03[3]), .C(n11528), .Z(n12697) );
  HS65_LL_NAND2X2 U14024 ( .A(n12697), .B(n13115), .Z(n12705) );
  HS65_LL_NAND2X2 U14025 ( .A(n11522), .B(n13104), .Z(n14575) );
  HS65_LL_NOR2X2 U14026 ( .A(sa03[6]), .B(n14575), .Z(n14903) );
  HS65_LL_NOR2X2 U14027 ( .A(sa03[0]), .B(sa03[3]), .Z(n14585) );
  HS65_LL_NAND2X2 U14028 ( .A(n14585), .B(n11528), .Z(n14925) );
  HS65_LL_NOR2X2 U14029 ( .A(n11544), .B(n14925), .Z(n14923) );
  HS65_LL_NOR2X2 U14030 ( .A(n11540), .B(n13119), .Z(n12711) );
  HS65_LL_NOR2X2 U14031 ( .A(n14923), .B(n12711), .Z(n11532) );
  HS65_LL_NOR3X1 U14032 ( .A(sa03[1]), .B(sa03[7]), .C(n12006), .Z(n13106) );
  HS65_LL_NAND2X2 U14033 ( .A(n12714), .B(n13106), .Z(n13781) );
  HS65_LL_NAND2X2 U14034 ( .A(n11532), .B(n13781), .Z(n12033) );
  HS65_LL_NOR4ABX2 U14035 ( .A(n11519), .B(n12705), .C(n14903), .D(n12033), 
        .Z(n14567) );
  HS65_LL_IVX2 U14036 ( .A(n14567), .Z(n12030) );
  HS65_LL_NOR3X1 U14037 ( .A(n15215), .B(n13099), .C(n12030), .Z(n11520) );
  HS65_LL_IVX2 U14038 ( .A(n12007), .Z(n12009) );
  HS65_LL_NAND2X2 U14039 ( .A(n11525), .B(n12009), .Z(n14905) );
  HS65_LL_IVX2 U14040 ( .A(n14594), .Z(n12713) );
  HS65_LL_NAND2X2 U14041 ( .A(n12697), .B(n12713), .Z(n14577) );
  HS65_LL_NAND3X2 U14042 ( .A(n11520), .B(n14905), .C(n14577), .Z(n11551) );
  HS65_LL_NOR2X2 U14043 ( .A(n14594), .B(n14925), .Z(n12715) );
  HS65_LL_NAND2X2 U14044 ( .A(n11521), .B(sa03[3]), .Z(n13120) );
  HS65_LL_OR2X4 U14045 ( .A(n13120), .B(sa03[5]), .Z(n14595) );
  HS65_LL_NOR2X2 U14046 ( .A(n12026), .B(n14595), .Z(n12702) );
  HS65_LL_NOR3X1 U14047 ( .A(sa03[5]), .B(n13120), .C(n13119), .Z(n13129) );
  HS65_LL_NOR2X2 U14048 ( .A(n12702), .B(n13129), .Z(n12728) );
  HS65_LL_IVX2 U14049 ( .A(n11548), .Z(n11536) );
  HS65_LL_NOR2X2 U14050 ( .A(n11536), .B(n12007), .Z(n14917) );
  HS65_LL_NOR2X2 U14051 ( .A(n12026), .B(n12007), .Z(n14573) );
  HS65_LL_NOR2X2 U14052 ( .A(n14917), .B(n14573), .Z(n12738) );
  HS65_LL_NOR2X2 U14053 ( .A(n11528), .B(n13120), .Z(n11545) );
  HS65_LL_NAND3X2 U14054 ( .A(sa03[7]), .B(n11545), .C(n11526), .Z(n14924) );
  HS65_LL_NOR2X2 U14055 ( .A(sa03[6]), .B(n14924), .Z(n14593) );
  HS65_LL_NAND2X2 U14056 ( .A(n11533), .B(n12713), .Z(n14581) );
  HS65_LL_IVX2 U14057 ( .A(n11545), .Z(n11534) );
  HS65_LL_NOR2X2 U14058 ( .A(n14574), .B(n11534), .Z(n15216) );
  HS65_LL_NAND2X2 U14059 ( .A(sa03[1]), .B(n15216), .Z(n12737) );
  HS65_LL_NAND2X2 U14060 ( .A(n14581), .B(n12737), .Z(n13795) );
  HS65_LL_NOR4ABX2 U14061 ( .A(n12728), .B(n12738), .C(n14593), .D(n13795), 
        .Z(n11523) );
  HS65_LL_IVX2 U14062 ( .A(n11522), .Z(n12726) );
  HS65_LL_NOR2X2 U14063 ( .A(sa03[6]), .B(n12726), .Z(n14584) );
  HS65_LL_NAND2X2 U14064 ( .A(n14584), .B(n12009), .Z(n15217) );
  HS65_LL_NAND2X2 U14065 ( .A(n13106), .B(n11545), .Z(n12036) );
  HS65_LL_NAND3X2 U14066 ( .A(n11523), .B(n15217), .C(n12036), .Z(n15208) );
  HS65_LL_NOR2X2 U14067 ( .A(n11534), .B(n14594), .Z(n15225) );
  HS65_LL_IVX2 U14068 ( .A(n12697), .Z(n12025) );
  HS65_LL_NOR2X2 U14069 ( .A(n12025), .B(n11536), .Z(n13108) );
  HS65_LL_NOR2X2 U14070 ( .A(n15225), .B(n13108), .Z(n13782) );
  HS65_LL_NAND2X2 U14071 ( .A(n12697), .B(n13105), .Z(n13785) );
  HS65_LL_NAND4ABX3 U14072 ( .A(n12715), .B(n15208), .C(n13782), .D(n13785), 
        .Z(n11524) );
  HS65_LL_NOR3X1 U14073 ( .A(sa03[5]), .B(n12022), .C(n14594), .Z(n12731) );
  HS65_LL_NOR3X1 U14074 ( .A(n11526), .B(n14574), .C(n14595), .Z(n12004) );
  HS65_LL_NOR2X2 U14075 ( .A(n12731), .B(n12004), .Z(n11531) );
  HS65_LL_NOR3X1 U14076 ( .A(sa03[5]), .B(n13120), .C(n12027), .Z(n14921) );
  HS65_LL_NOR2X2 U14077 ( .A(n11534), .B(n13119), .Z(n14611) );
  HS65_LL_NOR2X2 U14078 ( .A(n14921), .B(n14611), .Z(n12721) );
  HS65_LL_NAND4ABX3 U14079 ( .A(n11551), .B(n11524), .C(n11531), .D(n12721), 
        .Z(n11556) );
  HS65_LL_IVX2 U14080 ( .A(sa03[4]), .Z(n11543) );
  HS65_LL_NOR2X2 U14081 ( .A(sa03[2]), .B(n11543), .Z(n15238) );
  HS65_LL_NOR2X2 U14082 ( .A(n12027), .B(n14925), .Z(n14602) );
  HS65_LL_IVX2 U14083 ( .A(n15225), .Z(n13767) );
  HS65_LL_NAND2X2 U14084 ( .A(n11525), .B(n13104), .Z(n13772) );
  HS65_LL_NAND2X2 U14085 ( .A(n13767), .B(n13772), .Z(n11541) );
  HS65_LL_NAND2X2 U14086 ( .A(n14905), .B(n12720), .Z(n15199) );
  HS65_LL_NOR3X1 U14087 ( .A(sa03[6]), .B(n11526), .C(n14595), .Z(n13798) );
  HS65_LL_NOR3X1 U14088 ( .A(n11541), .B(n15199), .C(n13798), .Z(n11527) );
  HS65_LL_IVX2 U14089 ( .A(n12026), .Z(n12696) );
  HS65_LL_NAND2X2 U14090 ( .A(n12714), .B(n12696), .Z(n14918) );
  HS65_LL_NAND3AX3 U14091 ( .A(n14602), .B(n11527), .C(n14918), .Z(n15211) );
  HS65_LL_IVX2 U14092 ( .A(n12702), .Z(n12722) );
  HS65_LL_NAND2X2 U14093 ( .A(n12722), .B(n12737), .Z(n13103) );
  HS65_LL_NOR2X2 U14094 ( .A(n12007), .B(n13119), .Z(n14908) );
  HS65_LL_NOR3X1 U14095 ( .A(sa03[0]), .B(n11528), .C(n13119), .Z(n12021) );
  HS65_LL_IVX2 U14096 ( .A(n13106), .Z(n13790) );
  HS65_LL_NOR2X2 U14097 ( .A(n13790), .B(n11540), .Z(n13766) );
  HS65_LL_IVX2 U14098 ( .A(n13766), .Z(n11549) );
  HS65_LL_AOI12X2 U14099 ( .A(n12009), .B(n12695), .C(n14921), .Z(n11529) );
  HS65_LL_NAND4ABX3 U14100 ( .A(n14908), .B(n12021), .C(n11549), .D(n11529), 
        .Z(n11530) );
  HS65_LL_NOR3AX2 U14101 ( .A(n11531), .B(n13103), .C(n11530), .Z(n13788) );
  HS65_LL_OAI112X1 U14102 ( .A(n12022), .B(n11536), .C(n11532), .D(n13788), 
        .Z(n11535) );
  HS65_LL_NAND2X2 U14103 ( .A(n11533), .B(n14584), .Z(n13792) );
  HS65_LL_NOR2X2 U14104 ( .A(n12026), .B(n14925), .Z(n15205) );
  HS65_LL_NOR2AX3 U14105 ( .A(n13792), .B(n15205), .Z(n12040) );
  HS65_LL_IVX2 U14106 ( .A(n14584), .Z(n13111) );
  HS65_LL_NOR2X2 U14107 ( .A(n13111), .B(n14925), .Z(n12739) );
  HS65_LL_NOR2X2 U14108 ( .A(n13111), .B(n11534), .Z(n13094) );
  HS65_LL_NAND2X2 U14109 ( .A(n12714), .B(n13115), .Z(n15196) );
  HS65_LL_NAND2X2 U14110 ( .A(n12036), .B(n15196), .Z(n12010) );
  HS65_LL_NOR3X1 U14111 ( .A(n12739), .B(n13094), .C(n12010), .Z(n14570) );
  HS65_LL_NAND4ABX3 U14112 ( .A(n15211), .B(n11535), .C(n12040), .D(n14570), 
        .Z(n11555) );
  HS65_LL_NOR2X2 U14113 ( .A(sa03[2]), .B(sa03[4]), .Z(n15240) );
  HS65_LL_NOR2AX3 U14114 ( .A(n12714), .B(n13111), .Z(n13113) );
  HS65_LL_AND2X4 U14115 ( .A(n13104), .B(n12696), .Z(n13784) );
  HS65_LL_NOR2X2 U14116 ( .A(n12025), .B(n13111), .Z(n15227) );
  HS65_LL_NOR3X1 U14117 ( .A(n13113), .B(n13784), .C(n15227), .Z(n15214) );
  HS65_LL_NOR2X2 U14118 ( .A(n13120), .B(n12027), .Z(n11538) );
  HS65_LL_IVX2 U14119 ( .A(n13785), .Z(n14913) );
  HS65_LL_NOR2X2 U14120 ( .A(n11536), .B(n11540), .Z(n12028) );
  HS65_LL_NOR2X2 U14121 ( .A(n14913), .B(n12028), .Z(n13122) );
  HS65_LL_IVX2 U14122 ( .A(n13114), .Z(n12038) );
  HS65_LL_NOR3X1 U14123 ( .A(sa03[5]), .B(n12038), .C(n13790), .Z(n13780) );
  HS65_LL_NAND2X2 U14124 ( .A(n11549), .B(n15196), .Z(n12710) );
  HS65_LL_NOR4X4 U14125 ( .A(n13780), .B(n13108), .C(n13774), .D(n12710), .Z(
        n11537) );
  HS65_LL_NOR3X1 U14126 ( .A(sa03[1]), .B(n12006), .C(n14595), .Z(n15209) );
  HS65_LL_NAND2X2 U14127 ( .A(sa03[7]), .B(n15209), .Z(n12732) );
  HS65_LL_NAND3X2 U14128 ( .A(n13122), .B(n11537), .C(n12732), .Z(n14940) );
  HS65_LL_NOR3X1 U14129 ( .A(n11538), .B(n15215), .C(n14940), .Z(n11539) );
  HS65_LL_NAND3AX3 U14130 ( .A(n12711), .B(n15214), .C(n11539), .Z(n13098) );
  HS65_LL_NAND2X2 U14131 ( .A(n12714), .B(n11548), .Z(n12035) );
  HS65_LL_NAND2X2 U14132 ( .A(n12035), .B(n14577), .Z(n12013) );
  HS65_LL_NOR2X2 U14133 ( .A(n11540), .B(n12027), .Z(n14591) );
  HS65_LL_NOR3X1 U14134 ( .A(n14591), .B(n13129), .C(n12739), .Z(n12019) );
  HS65_LL_NOR2X2 U14135 ( .A(n12022), .B(n13790), .Z(n12017) );
  HS65_LL_IVX2 U14136 ( .A(n14923), .Z(n15206) );
  HS65_LL_NAND3AX3 U14137 ( .A(n11541), .B(n15206), .C(n14607), .Z(n13127) );
  HS65_LL_NOR4ABX2 U14138 ( .A(n12019), .B(n14905), .C(n12017), .D(n13127), 
        .Z(n11542) );
  HS65_LL_IVX2 U14139 ( .A(n12004), .Z(n12716) );
  HS65_LL_NAND4ABX3 U14140 ( .A(n13098), .B(n12013), .C(n11542), .D(n12716), 
        .Z(n11554) );
  HS65_LL_IVX2 U14141 ( .A(sa03[2]), .Z(n11552) );
  HS65_LL_NOR2X2 U14142 ( .A(n11552), .B(n11543), .Z(n15236) );
  HS65_LL_NOR2X2 U14143 ( .A(n11544), .B(n12025), .Z(n13095) );
  HS65_LL_IVX2 U14144 ( .A(n12035), .Z(n12703) );
  HS65_LL_NOR2X2 U14145 ( .A(n13095), .B(n12703), .Z(n14582) );
  HS65_LL_NOR2X2 U14146 ( .A(n12702), .B(n13780), .Z(n15229) );
  HS65_LL_NAND2X2 U14147 ( .A(n12696), .B(n11545), .Z(n12741) );
  HS65_LL_IVX2 U14148 ( .A(n14591), .Z(n12730) );
  HS65_LL_NAND2X2 U14149 ( .A(n12741), .B(n12730), .Z(n12694) );
  HS65_LL_NAND2X2 U14150 ( .A(n13105), .B(n12009), .Z(n14571) );
  HS65_LL_NAND2X2 U14151 ( .A(n13792), .B(n14571), .Z(n12736) );
  HS65_LL_NOR3X1 U14152 ( .A(n13129), .B(n12694), .C(n12736), .Z(n11546) );
  HS65_LL_NAND3X2 U14153 ( .A(n14582), .B(n15229), .C(n11546), .Z(n13118) );
  HS65_LL_IVX2 U14154 ( .A(n15216), .Z(n12037) );
  HS65_LL_NOR2X2 U14155 ( .A(sa03[1]), .B(n12037), .Z(n12018) );
  HS65_LL_NOR3X1 U14156 ( .A(n15225), .B(n12018), .C(n14602), .Z(n13097) );
  HS65_LL_IVX2 U14157 ( .A(n12739), .Z(n13107) );
  HS65_LL_NAND3X2 U14158 ( .A(n13097), .B(n13107), .C(n15217), .Z(n11547) );
  HS65_LL_NOR3X1 U14159 ( .A(n12715), .B(n14921), .C(n11547), .Z(n14937) );
  HS65_LL_IVX2 U14160 ( .A(n14925), .Z(n12712) );
  HS65_LL_NAND2X2 U14161 ( .A(n11548), .B(n12712), .Z(n15200) );
  HS65_LL_NAND2X2 U14162 ( .A(n14581), .B(n15200), .Z(n12699) );
  HS65_LL_NOR4ABX2 U14163 ( .A(n15214), .B(n11549), .C(n14917), .D(n12699), 
        .Z(n11550) );
  HS65_LL_NAND4ABX3 U14164 ( .A(n13118), .B(n11551), .C(n14937), .D(n11550), 
        .Z(n11553) );
  HS65_LL_NOR2X2 U14165 ( .A(sa03[4]), .B(n11552), .Z(n15234) );
  HS65_LL_MX41X4 U14166 ( .D0(n11556), .S0(n15238), .D1(n11555), .S1(n15240), 
        .D2(n11554), .S2(n15236), .D3(n11553), .S3(n15234), .Z(n15247) );
  HS65_LLS_XNOR2X3 U14167 ( .A(n15518), .B(n15247), .Z(n15674) );
  HS65_LL_OAI21X2 U14168 ( .A(n15674), .B(n11562), .C(n14808), .Z(n11561) );
  HS65_LL_IVX2 U14169 ( .A(text_in_r[10]), .Z(n11558) );
  HS65_LL_OAI212X3 U14170 ( .A(w3[10]), .B(text_in_r[10]), .C(n11559), .D(
        n11558), .E(ld_r), .Z(n11560) );
  HS65_LL_CBI4I1X3 U14171 ( .A(n11562), .B(n15674), .C(n11561), .D(n11560), 
        .Z(N52) );
  HS65_LL_IVX2 U14172 ( .A(w1[10]), .Z(n15035) );
  HS65_LL_MUXI21X2 U14173 ( .D0(w1[10]), .D1(n15035), .S0(n15451), .Z(n11563)
         );
  HS65_LLS_XOR3X2 U14174 ( .A(n14647), .B(n11563), .C(n15369), .Z(n11616) );
  HS65_LL_NOR2X2 U14175 ( .A(n11573), .B(n11564), .Z(n11571) );
  HS65_LL_OAI21X2 U14176 ( .A(n11602), .B(n11566), .C(n11565), .Z(n11567) );
  HS65_LL_NAND4ABX3 U14177 ( .A(n11798), .B(n11567), .C(n14423), .D(n11603), 
        .Z(n11568) );
  HS65_LL_NOR4ABX2 U14178 ( .A(n11571), .B(n11570), .C(n11569), .D(n11568), 
        .Z(n11612) );
  HS65_LL_NOR4ABX2 U14179 ( .A(n11575), .B(n11574), .C(n11573), .D(n11572), 
        .Z(n11589) );
  HS65_LL_NOR4ABX2 U14180 ( .A(n11589), .B(n14411), .C(n11577), .D(n11576), 
        .Z(n11578) );
  HS65_LL_NAND4ABX3 U14181 ( .A(n11581), .B(n11580), .C(n11579), .D(n11578), 
        .Z(n11591) );
  HS65_LL_NOR2AX3 U14182 ( .A(n11583), .B(n11582), .Z(n11596) );
  HS65_LL_NOR4ABX2 U14183 ( .A(n11596), .B(n11586), .C(n11585), .D(n11584), 
        .Z(n11588) );
  HS65_LL_AOI13X2 U14184 ( .A(n14444), .B(n11589), .C(n11588), .D(n11587), .Z(
        n11590) );
  HS65_LL_CBI4I6X2 U14185 ( .A(n11592), .B(n11591), .C(n14449), .D(n11590), 
        .Z(n11610) );
  HS65_LL_IVX2 U14186 ( .A(n11593), .Z(n11797) );
  HS65_LL_NOR4ABX2 U14187 ( .A(n11594), .B(n14411), .C(n11793), .D(n11797), 
        .Z(n11595) );
  HS65_LL_NAND4ABX3 U14188 ( .A(n11598), .B(n11597), .C(n11596), .D(n11595), 
        .Z(n14422) );
  HS65_LL_OAI112X1 U14189 ( .A(n11602), .B(n11601), .C(n11600), .D(n11599), 
        .Z(n11605) );
  HS65_LL_NAND4ABX3 U14190 ( .A(n11606), .B(n11605), .C(n11604), .D(n11603), 
        .Z(n11607) );
  HS65_LL_OAI13X1 U14191 ( .A(n14422), .B(n11608), .C(n11607), .D(n14453), .Z(
        n11609) );
  HS65_LL_OAI112X1 U14192 ( .A(n11612), .B(n11611), .C(n11610), .D(n11609), 
        .Z(n15133) );
  HS65_LLS_XNOR2X3 U14193 ( .A(n14854), .B(n15133), .Z(n14969) );
  HS65_LL_OAI21X2 U14194 ( .A(n14969), .B(n11616), .C(n14832), .Z(n11615) );
  HS65_LL_IVX2 U14195 ( .A(text_in_r[74]), .Z(n11613) );
  HS65_LL_OAI212X3 U14196 ( .A(w1[10]), .B(text_in_r[74]), .C(n15035), .D(
        n11613), .E(n15698), .Z(n11614) );
  HS65_LL_CBI4I1X3 U14197 ( .A(n11616), .B(n14969), .C(n11615), .D(n11614), 
        .Z(N180) );
  HS65_LL_MUX21I1X3 U14198 ( .D0(n11618), .D1(key[61]), .S0(n11617), .Z(
        \u0/N203 ) );
  HS65_LL_MUXI21X2 U14199 ( .D0(n15260), .D1(w0[17]), .S0(n14633), .Z(n11701)
         );
  HS65_LL_NAND4ABX3 U14200 ( .A(n13942), .B(n11619), .C(n13573), .D(n13943), 
        .Z(n11622) );
  HS65_LL_NOR4ABX2 U14201 ( .A(n12987), .B(n11620), .C(n12988), .D(n13597), 
        .Z(n11621) );
  HS65_LL_NAND4ABX3 U14202 ( .A(n11656), .B(n11622), .C(n13610), .D(n11621), 
        .Z(n11660) );
  HS65_LL_NOR2X2 U14203 ( .A(n11624), .B(n11623), .Z(n12424) );
  HS65_LL_NOR2X2 U14204 ( .A(n11625), .B(n13599), .Z(n12399) );
  HS65_LL_NAND4ABX3 U14205 ( .A(n11626), .B(n12424), .C(n12399), .D(n11636), 
        .Z(n11633) );
  HS65_LL_NAND4ABX3 U14206 ( .A(n13602), .B(n11628), .C(n11627), .D(n12410), 
        .Z(n11629) );
  HS65_LL_NOR4ABX2 U14207 ( .A(n11630), .B(n11635), .C(n12978), .D(n11629), 
        .Z(n12966) );
  HS65_LL_NAND4ABX3 U14208 ( .A(n11644), .B(n13970), .C(n12966), .D(n11631), 
        .Z(n11632) );
  HS65_LL_NOR2X2 U14209 ( .A(n12398), .B(n11641), .Z(n11651) );
  HS65_LL_NAND4ABX3 U14210 ( .A(n11633), .B(n11632), .C(n13610), .D(n11651), 
        .Z(n11659) );
  HS65_LL_NOR4ABX2 U14211 ( .A(n11636), .B(n11635), .C(n13003), .D(n11634), 
        .Z(n13607) );
  HS65_LL_NOR4ABX2 U14212 ( .A(n13607), .B(n11638), .C(n11637), .D(n13602), 
        .Z(n11640) );
  HS65_LL_NAND4ABX3 U14213 ( .A(n11641), .B(n12968), .C(n11640), .D(n11639), 
        .Z(n13959) );
  HS65_LL_NOR2X2 U14214 ( .A(n13599), .B(n12981), .Z(n13949) );
  HS65_LL_NOR2X2 U14215 ( .A(n13571), .B(n11642), .Z(n12992) );
  HS65_LL_NAND2AX4 U14216 ( .A(n11644), .B(n11643), .Z(n12397) );
  HS65_LL_NAND2X2 U14217 ( .A(n11645), .B(n12405), .Z(n13587) );
  HS65_LL_NOR4ABX2 U14218 ( .A(n13949), .B(n12992), .C(n12397), .D(n13587), 
        .Z(n11647) );
  HS65_LL_NAND4ABX3 U14219 ( .A(n13959), .B(n11648), .C(n11647), .D(n11646), 
        .Z(n11658) );
  HS65_LL_NOR2X2 U14220 ( .A(n11650), .B(n11649), .Z(n12413) );
  HS65_LL_NAND4ABX3 U14221 ( .A(n12413), .B(n13598), .C(n11651), .D(n13566), 
        .Z(n11655) );
  HS65_LL_NOR4ABX2 U14222 ( .A(n13573), .B(n13968), .C(n11652), .D(n13971), 
        .Z(n11653) );
  HS65_LL_NAND4ABX3 U14223 ( .A(n11656), .B(n11655), .C(n11654), .D(n11653), 
        .Z(n11657) );
  HS65_LL_MX41X4 U14224 ( .D0(n11660), .S0(n13961), .D1(n11659), .S1(n13972), 
        .D2(n11658), .S2(n13614), .D3(n11657), .S3(n13981), .Z(n15261) );
  HS65_LL_IVX2 U14225 ( .A(n15261), .Z(n15262) );
  HS65_LL_MUXI21X2 U14226 ( .D0(n15262), .D1(n15261), .S0(n15552), .Z(n11700)
         );
  HS65_LL_IVX2 U14227 ( .A(n15251), .Z(n15252) );
  HS65_LL_NOR4ABX2 U14228 ( .A(n12495), .B(n11661), .C(n12439), .D(n12926), 
        .Z(n11662) );
  HS65_LL_NAND4ABX3 U14229 ( .A(n12514), .B(n11664), .C(n11663), .D(n11662), 
        .Z(n11699) );
  HS65_LL_AND2X4 U14230 ( .A(n12527), .B(n11665), .Z(n12461) );
  HS65_LL_AOI13X2 U14231 ( .A(n11745), .B(sa22[7]), .C(n11667), .D(n11666), 
        .Z(n11676) );
  HS65_LL_IVX2 U14232 ( .A(n12492), .Z(n11668) );
  HS65_LL_NAND4ABX3 U14233 ( .A(n11671), .B(n11670), .C(n11669), .D(n11668), 
        .Z(n11757) );
  HS65_LL_NOR4ABX2 U14234 ( .A(n11672), .B(n12454), .C(n12476), .D(n12505), 
        .Z(n11673) );
  HS65_LL_OAI21X2 U14235 ( .A(n11675), .B(n11674), .C(n11673), .Z(n11754) );
  HS65_LL_NOR4ABX2 U14236 ( .A(n12461), .B(n11676), .C(n11757), .D(n11754), 
        .Z(n11677) );
  HS65_LL_NAND2X2 U14237 ( .A(n11678), .B(n11677), .Z(n11698) );
  HS65_LL_NAND2X2 U14238 ( .A(n12480), .B(n11679), .Z(n11681) );
  HS65_LL_NAND4ABX3 U14239 ( .A(n12446), .B(n11681), .C(n11680), .D(n12443), 
        .Z(n11687) );
  HS65_LL_NAND3X2 U14240 ( .A(n11684), .B(n11683), .C(n11682), .Z(n11685) );
  HS65_LL_NOR3X1 U14241 ( .A(n11689), .B(n12460), .C(n11685), .Z(n12518) );
  HS65_LL_NAND4ABX3 U14242 ( .A(n12519), .B(n11687), .C(n12518), .D(n11686), 
        .Z(n11697) );
  HS65_LL_IVX2 U14243 ( .A(n12526), .Z(n11752) );
  HS65_LL_NOR4ABX2 U14244 ( .A(n11690), .B(n11752), .C(n11689), .D(n11688), 
        .Z(n11691) );
  HS65_LL_NOR4ABX2 U14245 ( .A(n11692), .B(n11691), .C(n12485), .D(n12936), 
        .Z(n11693) );
  HS65_LL_NAND3X2 U14246 ( .A(n11695), .B(n11694), .C(n11693), .Z(n11696) );
  HS65_LL_MX41X4 U14247 ( .D0(n11699), .S0(n12540), .D1(n11698), .S1(n12951), 
        .D2(n11697), .S2(n12943), .D3(n11696), .S3(n12945), .Z(n15345) );
  HS65_LL_MUXI21X2 U14248 ( .D0(n15251), .D1(n15252), .S0(n15345), .Z(n13855)
         );
  HS65_LLS_XOR3X2 U14249 ( .A(n11701), .B(n11700), .C(n13855), .Z(n11772) );
  HS65_LL_NAND3X2 U14250 ( .A(n11703), .B(n11702), .C(n13527), .Z(n13510) );
  HS65_LL_NOR3X1 U14251 ( .A(n13541), .B(n12603), .C(n13510), .Z(n14042) );
  HS65_LL_NOR4ABX2 U14252 ( .A(n11704), .B(n13539), .C(n11715), .D(n13650), 
        .Z(n11705) );
  HS65_LL_NAND4ABX3 U14253 ( .A(n14069), .B(n11706), .C(n14042), .D(n11705), 
        .Z(n11735) );
  HS65_LL_NAND2X2 U14254 ( .A(n13544), .B(n11707), .Z(n14043) );
  HS65_LL_IVX2 U14255 ( .A(n11715), .Z(n13534) );
  HS65_LL_NAND2X2 U14256 ( .A(n13534), .B(n13506), .Z(n13628) );
  HS65_LL_NOR4ABX2 U14257 ( .A(n11709), .B(n11708), .C(n13639), .D(n13628), 
        .Z(n11710) );
  HS65_LL_NAND4ABX3 U14258 ( .A(n13524), .B(n14043), .C(n11711), .D(n11710), 
        .Z(n11734) );
  HS65_LL_NOR2X2 U14259 ( .A(n11712), .B(n13543), .Z(n13622) );
  HS65_LL_NOR4ABX2 U14260 ( .A(n13622), .B(n11714), .C(n14030), .D(n11713), 
        .Z(n13514) );
  HS65_LL_NOR2X2 U14261 ( .A(n11715), .B(n14033), .Z(n14063) );
  HS65_LL_NOR4ABX2 U14262 ( .A(n13538), .B(n14063), .C(n11717), .D(n11716), 
        .Z(n11718) );
  HS65_LL_NAND4ABX3 U14263 ( .A(n11731), .B(n11719), .C(n13514), .D(n11718), 
        .Z(n11733) );
  HS65_LL_OAI112X1 U14264 ( .A(n11722), .B(n11721), .C(n11720), .D(n13641), 
        .Z(n12605) );
  HS65_LL_NOR2X2 U14265 ( .A(n11723), .B(n13553), .Z(n13520) );
  HS65_LL_OAI112X1 U14266 ( .A(n13559), .B(n11725), .C(n11724), .D(n13520), 
        .Z(n11726) );
  HS65_LL_NOR4ABX2 U14267 ( .A(n13621), .B(n12600), .C(n12605), .D(n11726), 
        .Z(n13653) );
  HS65_LL_AND2X4 U14268 ( .A(n11727), .B(n13548), .Z(n14045) );
  HS65_LL_NOR4ABX2 U14269 ( .A(n14045), .B(n12622), .C(n12621), .D(n11728), 
        .Z(n11729) );
  HS65_LL_NAND4ABX3 U14270 ( .A(n11731), .B(n11730), .C(n13653), .D(n11729), 
        .Z(n11732) );
  HS65_LL_MX41X4 U14271 ( .D0(n11735), .S0(n13659), .D1(n11734), .S1(n13657), 
        .D2(n11733), .S2(n14067), .D3(n11732), .S3(n14075), .Z(n15441) );
  HS65_LL_IVX2 U14272 ( .A(n15441), .Z(n15442) );
  HS65_LL_NOR3X1 U14273 ( .A(n11751), .B(n11761), .C(n11736), .Z(n12914) );
  HS65_LL_NOR4ABX2 U14274 ( .A(n12914), .B(n11739), .C(n11738), .D(n11737), 
        .Z(n11740) );
  HS65_LL_NAND4ABX3 U14275 ( .A(n11754), .B(n11742), .C(n11741), .D(n11740), 
        .Z(n11768) );
  HS65_LL_NOR2X2 U14276 ( .A(n11743), .B(n12530), .Z(n12932) );
  HS65_LL_AOI12X2 U14277 ( .A(n11746), .B(n11745), .C(n11744), .Z(n12475) );
  HS65_LL_NAND4ABX3 U14278 ( .A(n11747), .B(n12440), .C(n12466), .D(n12475), 
        .Z(n11748) );
  HS65_LL_NOR4ABX2 U14279 ( .A(n12467), .B(n12461), .C(n11749), .D(n11748), 
        .Z(n12456) );
  HS65_LL_NOR4ABX2 U14280 ( .A(n12456), .B(n11752), .C(n11751), .D(n11750), 
        .Z(n11753) );
  HS65_LL_NAND4ABX3 U14281 ( .A(n11754), .B(n12468), .C(n12932), .D(n11753), 
        .Z(n11767) );
  HS65_LL_NOR3X1 U14282 ( .A(n12498), .B(n11756), .C(n11755), .Z(n11758) );
  HS65_LL_NOR4ABX2 U14283 ( .A(n12518), .B(n11758), .C(n11761), .D(n11757), 
        .Z(n11759) );
  HS65_LL_NAND3X2 U14284 ( .A(n12920), .B(n12909), .C(n11759), .Z(n11766) );
  HS65_LL_NOR2X2 U14285 ( .A(n11761), .B(n11760), .Z(n12463) );
  HS65_LL_NOR4ABX2 U14286 ( .A(n12463), .B(n12443), .C(n12526), .D(n12451), 
        .Z(n11762) );
  HS65_LL_NAND4ABX3 U14287 ( .A(n11764), .B(n12519), .C(n11763), .D(n11762), 
        .Z(n11765) );
  HS65_LL_MX41X4 U14288 ( .D0(n11768), .S0(n12540), .D1(n11767), .S1(n12951), 
        .D2(n11766), .S2(n12943), .D3(n11765), .S3(n12945), .Z(n15355) );
  HS65_LL_MUXI21X2 U14289 ( .D0(n15442), .D1(n15441), .S0(n15355), .Z(n15536)
         );
  HS65_LL_OAI21X2 U14290 ( .A(n15536), .B(n11772), .C(n14808), .Z(n11771) );
  HS65_LL_IVX2 U14291 ( .A(text_in_r[113]), .Z(n11769) );
  HS65_LL_OAI212X3 U14292 ( .A(w0[17]), .B(text_in_r[113]), .C(n15260), .D(
        n11769), .E(n15698), .Z(n11770) );
  HS65_LL_CBI4I1X3 U14293 ( .A(n11772), .B(n15536), .C(n11771), .D(n11770), 
        .Z(N259) );
  HS65_LL_NOR2X2 U14294 ( .A(sa01[7]), .B(n11773), .Z(n11775) );
  HS65_LL_AOI112X2 U14295 ( .A(n11776), .B(n11775), .C(n11774), .D(n14421), 
        .Z(n11777) );
  HS65_LL_NAND4ABX3 U14296 ( .A(n11779), .B(n14415), .C(n11778), .D(n11777), 
        .Z(n11813) );
  HS65_LL_NAND4ABX3 U14297 ( .A(n11783), .B(n11782), .C(n11781), .D(n11780), 
        .Z(n11786) );
  HS65_LL_NAND4ABX3 U14298 ( .A(n11787), .B(n11786), .C(n11785), .D(n11784), 
        .Z(n11812) );
  HS65_LL_AND2X4 U14299 ( .A(n11789), .B(n11788), .Z(n14418) );
  HS65_LL_NOR2X2 U14300 ( .A(n14442), .B(n11790), .Z(n11791) );
  HS65_LL_NAND4ABX3 U14301 ( .A(n11794), .B(n11793), .C(n11792), .D(n11791), 
        .Z(n11795) );
  HS65_LL_NOR4ABX2 U14302 ( .A(n11796), .B(n14418), .C(n11804), .D(n11795), 
        .Z(n14429) );
  HS65_LL_NOR4ABX2 U14303 ( .A(n11799), .B(n14408), .C(n11798), .D(n11797), 
        .Z(n11800) );
  HS65_LL_NAND4ABX3 U14304 ( .A(n11809), .B(n11801), .C(n14429), .D(n11800), 
        .Z(n11811) );
  HS65_LL_NAND4ABX3 U14305 ( .A(n11805), .B(n11804), .C(n11803), .D(n11802), 
        .Z(n11808) );
  HS65_LL_NAND4ABX3 U14306 ( .A(n11809), .B(n11808), .C(n11807), .D(n11806), 
        .Z(n11810) );
  HS65_LL_MX41X4 U14307 ( .D0(n11813), .S0(n14453), .D1(n11812), .S1(n14451), 
        .D2(n11811), .S2(n14449), .D3(n11810), .S3(n14447), .Z(n15135) );
  HS65_LLS_XOR2X3 U14308 ( .A(n15135), .B(n15451), .Z(n14961) );
  HS65_LL_IVX2 U14309 ( .A(n15275), .Z(n15276) );
  HS65_LL_IVX2 U14310 ( .A(n11814), .Z(n12223) );
  HS65_LL_NAND2X2 U14311 ( .A(n14330), .B(n14302), .Z(n11839) );
  HS65_LL_NAND2X2 U14312 ( .A(n11816), .B(n11815), .Z(n12211) );
  HS65_LL_NOR3X1 U14313 ( .A(n11817), .B(n11871), .C(n12211), .Z(n14311) );
  HS65_LL_NOR4ABX2 U14314 ( .A(n11819), .B(n11833), .C(n11818), .D(n13421), 
        .Z(n11820) );
  HS65_LL_NAND3X2 U14315 ( .A(n11820), .B(n12196), .C(n13423), .Z(n11821) );
  HS65_LL_NOR3X1 U14316 ( .A(n12205), .B(n11854), .C(n11821), .Z(n14293) );
  HS65_LL_NOR4ABX2 U14317 ( .A(n14293), .B(n11840), .C(n13414), .D(n11822), 
        .Z(n11823) );
  HS65_LL_NAND4ABX3 U14318 ( .A(n12223), .B(n11839), .C(n14311), .D(n11823), 
        .Z(n11852) );
  HS65_LL_NOR4ABX2 U14319 ( .A(n11833), .B(n11825), .C(n12200), .D(n11824), 
        .Z(n11897) );
  HS65_LL_NOR4ABX2 U14320 ( .A(n11829), .B(n11828), .C(n11827), .D(n11826), 
        .Z(n11830) );
  HS65_LL_NAND4ABX3 U14321 ( .A(n12223), .B(n11831), .C(n11897), .D(n11830), 
        .Z(n11851) );
  HS65_LL_NOR2X2 U14322 ( .A(n13429), .B(n11832), .Z(n13454) );
  HS65_LL_NAND2X2 U14323 ( .A(n11834), .B(n11833), .Z(n11886) );
  HS65_LL_NOR4ABX2 U14324 ( .A(n13454), .B(n11836), .C(n11886), .D(n11835), 
        .Z(n11837) );
  HS65_LL_NAND4ABX3 U14325 ( .A(n13438), .B(n11839), .C(n11838), .D(n11837), 
        .Z(n11850) );
  HS65_LL_NAND3X2 U14326 ( .A(n11842), .B(n11841), .C(n11840), .Z(n12212) );
  HS65_LL_NOR4ABX2 U14327 ( .A(n11875), .B(n11844), .C(n12212), .D(n11843), 
        .Z(n11846) );
  HS65_LL_NAND4ABX3 U14328 ( .A(n11848), .B(n11847), .C(n11846), .D(n11845), 
        .Z(n11849) );
  HS65_LL_MX41X4 U14329 ( .D0(n11852), .S0(n14337), .D1(n11851), .S1(n14339), 
        .D2(n11850), .S2(n14335), .D3(n11849), .S3(n14333), .Z(n15371) );
  HS65_LL_MUXI21X2 U14330 ( .D0(n15276), .D1(n15275), .S0(n15371), .Z(n14972)
         );
  HS65_LL_IVX2 U14331 ( .A(w1[17]), .Z(n15274) );
  HS65_LL_MUXI21X2 U14332 ( .D0(n15274), .D1(w1[17]), .S0(n15369), .Z(n11853)
         );
  HS65_LLS_XOR3X2 U14333 ( .A(n14961), .B(n14972), .C(n11853), .Z(n11901) );
  HS65_LL_NOR3X1 U14334 ( .A(n13428), .B(n11884), .C(n11854), .Z(n14315) );
  HS65_LL_AOI112X2 U14335 ( .A(n11856), .B(sa23[7]), .C(n13433), .D(n11855), 
        .Z(n11859) );
  HS65_LL_NOR4ABX2 U14336 ( .A(n14315), .B(n11859), .C(n11858), .D(n11857), 
        .Z(n11896) );
  HS65_LL_NAND3X2 U14337 ( .A(n14330), .B(n13453), .C(n11860), .Z(n11861) );
  HS65_LL_NOR3X1 U14338 ( .A(n14295), .B(n11862), .C(n11861), .Z(n14324) );
  HS65_LL_NOR2X2 U14339 ( .A(n11864), .B(n11863), .Z(n11865) );
  HS65_LL_NOR4ABX2 U14340 ( .A(n11867), .B(n14297), .C(n11866), .D(n11865), 
        .Z(n11868) );
  HS65_LL_NOR4ABX2 U14341 ( .A(n11876), .B(n11868), .C(n12205), .D(n13456), 
        .Z(n11869) );
  HS65_LL_NAND4ABX3 U14342 ( .A(n11871), .B(n11870), .C(n14324), .D(n11869), 
        .Z(n11894) );
  HS65_LL_NAND3X2 U14343 ( .A(n11873), .B(n14320), .C(n11872), .Z(n12219) );
  HS65_LL_NAND3X2 U14344 ( .A(n11876), .B(n11875), .C(n11874), .Z(n11877) );
  HS65_LL_NOR3X1 U14345 ( .A(n13433), .B(n12219), .C(n11877), .Z(n14329) );
  HS65_LL_NOR4ABX2 U14346 ( .A(n14315), .B(n13423), .C(n11879), .D(n11878), 
        .Z(n11881) );
  HS65_LL_AOI13X2 U14347 ( .A(n11882), .B(n14329), .C(n11881), .D(n11880), .Z(
        n11893) );
  HS65_LL_NOR2X2 U14348 ( .A(n11884), .B(n11883), .Z(n13425) );
  HS65_LL_NOR4ABX2 U14349 ( .A(n11887), .B(n13425), .C(n11886), .D(n11885), 
        .Z(n11889) );
  HS65_LL_AOI13X2 U14350 ( .A(n11891), .B(n11890), .C(n11889), .D(n11888), .Z(
        n11892) );
  HS65_LL_AOI112X2 U14351 ( .A(n14337), .B(n11894), .C(n11893), .D(n11892), 
        .Z(n11895) );
  HS65_LL_CBI4I1X3 U14352 ( .A(n11897), .B(n11896), .C(n12229), .D(n11895), 
        .Z(n15357) );
  HS65_LLS_XNOR2X3 U14353 ( .A(n15264), .B(n15357), .Z(n14964) );
  HS65_LL_OAI21X2 U14354 ( .A(n14964), .B(n11901), .C(n14832), .Z(n11900) );
  HS65_LL_IVX2 U14355 ( .A(text_in_r[81]), .Z(n11898) );
  HS65_LL_OAI212X3 U14356 ( .A(w1[17]), .B(text_in_r[81]), .C(n15274), .D(
        n11898), .E(n15545), .Z(n11899) );
  HS65_LL_CBI4I1X3 U14357 ( .A(n11901), .B(n14964), .C(n11900), .D(n11899), 
        .Z(N195) );
  HS65_LL_OAI21X2 U14358 ( .A(w1[31]), .B(text_in_r[95]), .C(n15698), .Z(
        n11906) );
  HS65_LL_IVX2 U14359 ( .A(n15357), .Z(n15358) );
  HS65_LL_MUXI21X2 U14360 ( .D0(n15357), .D1(n15358), .S0(n15443), .Z(n11902)
         );
  HS65_LL_NOR2AX3 U14361 ( .A(n11902), .B(n15698), .Z(n14858) );
  HS65_LL_NOR2X2 U14362 ( .A(n14822), .B(n11902), .Z(n14857) );
  HS65_LL_IVX2 U14363 ( .A(w1[31]), .Z(n15091) );
  HS65_LL_IVX2 U14364 ( .A(n15266), .Z(n15265) );
  HS65_LL_MUXI21X2 U14365 ( .D0(n15266), .D1(n15265), .S0(n15125), .Z(n14949)
         );
  HS65_LL_MUXI21X2 U14366 ( .D0(w1[31]), .D1(n15091), .S0(n14949), .Z(n11903)
         );
  HS65_LL_MUXI21X2 U14367 ( .D0(n15263), .D1(n15264), .S0(n11903), .Z(n11904)
         );
  HS65_LL_MUXI21X2 U14368 ( .D0(n14858), .D1(n14857), .S0(n11904), .Z(n11905)
         );
  HS65_LL_CBI4I1X3 U14369 ( .A(text_in_r[95]), .B(w1[31]), .C(n11906), .D(
        n11905), .Z(N217) );
  HS65_LL_IVX2 U14370 ( .A(n14166), .Z(n13224) );
  HS65_LL_NOR2X2 U14371 ( .A(n13239), .B(n13224), .Z(n12678) );
  HS65_LL_NAND2X2 U14372 ( .A(n12678), .B(n12656), .Z(n11930) );
  HS65_LL_IVX2 U14373 ( .A(n13231), .Z(n12665) );
  HS65_LL_IVX2 U14374 ( .A(n13817), .Z(n14242) );
  HS65_LL_NOR2X2 U14375 ( .A(n12683), .B(n14242), .Z(n12655) );
  HS65_LL_NAND3X2 U14376 ( .A(n12655), .B(n14173), .C(n11907), .Z(n11908) );
  HS65_LL_NOR3X1 U14377 ( .A(n11943), .B(n12665), .C(n11908), .Z(n13877) );
  HS65_LL_NAND4ABX3 U14378 ( .A(n14144), .B(n11930), .C(n13877), .D(n11940), 
        .Z(n11909) );
  HS65_LL_AOI12X2 U14379 ( .A(n11911), .B(n11910), .C(n11909), .Z(n14262) );
  HS65_LL_NAND2X2 U14380 ( .A(n12664), .B(n13228), .Z(n11912) );
  HS65_LL_NOR4ABX2 U14381 ( .A(n13220), .B(n12650), .C(n11913), .D(n11912), 
        .Z(n11920) );
  HS65_LL_IVX2 U14382 ( .A(n13860), .Z(n14243) );
  HS65_LL_NAND2X2 U14383 ( .A(n14243), .B(n11927), .Z(n11949) );
  HS65_LL_NOR4ABX2 U14384 ( .A(n11914), .B(n11937), .C(n13820), .D(n11949), 
        .Z(n11919) );
  HS65_LL_NAND2X2 U14385 ( .A(n13209), .B(n14240), .Z(n12660) );
  HS65_LL_NAND2AX4 U14386 ( .A(n13234), .B(n13235), .Z(n11918) );
  HS65_LL_NOR2X2 U14387 ( .A(n13839), .B(n13840), .Z(n11917) );
  HS65_LL_NOR4ABX2 U14388 ( .A(n12680), .B(n13229), .C(n13213), .D(n11915), 
        .Z(n11916) );
  HS65_LL_NAND4ABX3 U14389 ( .A(n12689), .B(n11918), .C(n11917), .D(n11916), 
        .Z(n14168) );
  HS65_LL_NOR4ABX2 U14390 ( .A(n11920), .B(n11919), .C(n12660), .D(n14168), 
        .Z(n11957) );
  HS65_LL_IVX2 U14391 ( .A(n14285), .Z(n11956) );
  HS65_LL_IVX2 U14392 ( .A(n13236), .Z(n14160) );
  HS65_LL_IVX2 U14393 ( .A(n11921), .Z(n13868) );
  HS65_LL_NAND2X2 U14394 ( .A(n13868), .B(n12647), .Z(n11947) );
  HS65_LL_NOR2X2 U14395 ( .A(n11942), .B(n11922), .Z(n14162) );
  HS65_LL_NAND2X2 U14396 ( .A(n14266), .B(n11923), .Z(n13841) );
  HS65_LL_NAND2X2 U14397 ( .A(n13841), .B(n12650), .Z(n13208) );
  HS65_LL_NOR3X1 U14398 ( .A(n14162), .B(n11924), .C(n13208), .Z(n11925) );
  HS65_LL_NAND4ABX3 U14399 ( .A(n14160), .B(n11947), .C(n11925), .D(n14257), 
        .Z(n13882) );
  HS65_LL_NAND2X2 U14400 ( .A(n11926), .B(n14151), .Z(n14253) );
  HS65_LL_NAND2X2 U14401 ( .A(n14253), .B(n11927), .Z(n12654) );
  HS65_LL_NOR2X2 U14402 ( .A(n13820), .B(n12654), .Z(n13869) );
  HS65_LL_NAND3X2 U14403 ( .A(n13221), .B(n13824), .C(n13818), .Z(n14183) );
  HS65_LL_NOR4ABX2 U14404 ( .A(n11934), .B(n13229), .C(n11928), .D(n14183), 
        .Z(n11929) );
  HS65_LL_NAND4ABX3 U14405 ( .A(n13882), .B(n11930), .C(n13869), .D(n11929), 
        .Z(n11954) );
  HS65_LL_NAND2X2 U14406 ( .A(n14243), .B(n14253), .Z(n14273) );
  HS65_LL_NAND2X2 U14407 ( .A(n13818), .B(n13235), .Z(n14153) );
  HS65_LL_NOR4X4 U14408 ( .A(n11932), .B(n14144), .C(n14278), .D(n11931), .Z(
        n13836) );
  HS65_LL_NAND4ABX3 U14409 ( .A(n13233), .B(n14153), .C(n13836), .D(n13206), 
        .Z(n11933) );
  HS65_LL_NOR4ABX2 U14410 ( .A(n11935), .B(n11934), .C(n14273), .D(n11933), 
        .Z(n11952) );
  HS65_LL_IVX2 U14411 ( .A(n14283), .Z(n11951) );
  HS65_LL_NAND2X2 U14412 ( .A(n13229), .B(n12651), .Z(n12673) );
  HS65_LL_NAND2X2 U14413 ( .A(n11936), .B(n13828), .Z(n14145) );
  HS65_LL_NOR4ABX2 U14414 ( .A(n14157), .B(n11937), .C(n14162), .D(n14145), 
        .Z(n13865) );
  HS65_LL_IVX2 U14415 ( .A(n14252), .Z(n13232) );
  HS65_LL_NAND2X2 U14416 ( .A(n12670), .B(n11938), .Z(n14150) );
  HS65_LL_NAND4ABX3 U14417 ( .A(n13232), .B(n14150), .C(n12664), .D(n13228), 
        .Z(n11939) );
  HS65_LL_NOR4ABX2 U14418 ( .A(n13865), .B(n11940), .C(n13239), .D(n11939), 
        .Z(n13823) );
  HS65_LL_IVX2 U14419 ( .A(n13200), .Z(n11944) );
  HS65_LL_NOR2X2 U14420 ( .A(n11942), .B(n11941), .Z(n14161) );
  HS65_LL_NOR2X2 U14421 ( .A(n11943), .B(n13233), .Z(n12682) );
  HS65_LL_NAND2AX4 U14422 ( .A(n14161), .B(n12682), .Z(n13890) );
  HS65_LL_NOR4ABX2 U14423 ( .A(n13823), .B(n11944), .C(n14144), .D(n13890), 
        .Z(n11946) );
  HS65_LL_NAND4ABX3 U14424 ( .A(n14256), .B(n11947), .C(n11946), .D(n11945), 
        .Z(n11948) );
  HS65_LL_OAI13X1 U14425 ( .A(n11949), .B(n12673), .C(n11948), .D(n14279), .Z(
        n11950) );
  HS65_LL_CBI4I1X3 U14426 ( .A(n14175), .B(n11952), .C(n11951), .D(n11950), 
        .Z(n11953) );
  HS65_LL_CBI4I6X2 U14427 ( .A(n12668), .B(n11954), .C(n14281), .D(n11953), 
        .Z(n11955) );
  HS65_LL_CBI4I1X3 U14428 ( .A(n14262), .B(n11957), .C(n11956), .D(n11955), 
        .Z(n15677) );
  HS65_LL_IVX2 U14429 ( .A(n15677), .Z(n15726) );
  HS65_LL_NAND2X2 U14430 ( .A(n11958), .B(n11986), .Z(n14873) );
  HS65_LL_NAND2X2 U14431 ( .A(n14873), .B(n13151), .Z(n11988) );
  HS65_LL_NOR4ABX2 U14432 ( .A(n11959), .B(n14215), .C(n14889), .D(n11988), 
        .Z(n12803) );
  HS65_LL_IVX2 U14433 ( .A(n11996), .Z(n12783) );
  HS65_LL_NOR2AX3 U14434 ( .A(n12103), .B(n12781), .Z(n12787) );
  HS65_LL_NAND3X2 U14435 ( .A(n11961), .B(n11989), .C(n11960), .Z(n12779) );
  HS65_LL_AOI112X2 U14436 ( .A(n12783), .B(n11962), .C(n12787), .D(n12779), 
        .Z(n11971) );
  HS65_LL_NOR3AX2 U14437 ( .A(n12132), .B(n11964), .C(n11963), .Z(n11976) );
  HS65_LL_NOR3X1 U14438 ( .A(n13903), .B(n11976), .C(n12784), .Z(n12762) );
  HS65_LL_IVX2 U14439 ( .A(n12750), .Z(n12796) );
  HS65_LL_NOR2X2 U14440 ( .A(n11966), .B(n11965), .Z(n12791) );
  HS65_LL_IVX2 U14441 ( .A(n12791), .Z(n11987) );
  HS65_LL_NAND2X2 U14442 ( .A(n11987), .B(n12128), .Z(n13149) );
  HS65_LL_NOR4ABX2 U14443 ( .A(n12796), .B(n13916), .C(n14864), .D(n13149), 
        .Z(n12118) );
  HS65_LL_IVX2 U14444 ( .A(n12131), .Z(n12752) );
  HS65_LL_NOR2X2 U14445 ( .A(n12114), .B(n12780), .Z(n11967) );
  HS65_LL_NAND4ABX3 U14446 ( .A(n13905), .B(n12108), .C(n11968), .D(n11967), 
        .Z(n11969) );
  HS65_LL_NOR4ABX2 U14447 ( .A(n12762), .B(n12118), .C(n12752), .D(n11969), 
        .Z(n11970) );
  HS65_LL_NAND3X2 U14448 ( .A(n12803), .B(n11971), .C(n11970), .Z(n12003) );
  HS65_LL_NAND3X2 U14449 ( .A(n11972), .B(n12105), .C(n14188), .Z(n11983) );
  HS65_LL_NOR2X2 U14450 ( .A(n13899), .B(n13156), .Z(n11973) );
  HS65_LL_NOR4ABX2 U14451 ( .A(n11973), .B(n11995), .C(n12795), .D(n13906), 
        .Z(n11974) );
  HS65_LL_NOR4ABX2 U14452 ( .A(n11974), .B(n12104), .C(n13904), .D(n12121), 
        .Z(n14228) );
  HS65_LL_IVX2 U14453 ( .A(n13164), .Z(n11993) );
  HS65_LL_NOR4ABX2 U14454 ( .A(n14873), .B(n11993), .C(n12114), .D(n12780), 
        .Z(n14887) );
  HS65_LL_NAND4ABX3 U14455 ( .A(n12134), .B(n11975), .C(n14228), .D(n14887), 
        .Z(n11982) );
  HS65_LL_NOR3X1 U14456 ( .A(n12101), .B(n14219), .C(n13149), .Z(n12773) );
  HS65_LL_NOR3X1 U14457 ( .A(n14872), .B(n12799), .C(n11992), .Z(n11977) );
  HS65_LL_NOR4ABX2 U14458 ( .A(n11977), .B(n12770), .C(n12758), .D(n11976), 
        .Z(n13928) );
  HS65_LL_CBI4I1X3 U14459 ( .A(n11980), .B(n11979), .C(n11978), .D(n12769), 
        .Z(n11981) );
  HS65_LL_NOR3AX2 U14460 ( .A(n13928), .B(n11998), .C(n11981), .Z(n14194) );
  HS65_LL_NAND4ABX3 U14461 ( .A(n11983), .B(n11982), .C(n12773), .D(n14194), 
        .Z(n12002) );
  HS65_LL_NAND2X2 U14462 ( .A(n11984), .B(n14188), .Z(n12113) );
  HS65_LL_IVX2 U14463 ( .A(n11995), .Z(n14871) );
  HS65_LL_NOR2X2 U14464 ( .A(n14863), .B(n14871), .Z(n11991) );
  HS65_LL_NAND2X2 U14465 ( .A(n12105), .B(n14220), .Z(n12778) );
  HS65_LL_NAND2X2 U14466 ( .A(n12119), .B(n12788), .Z(n14222) );
  HS65_LL_OAI21X2 U14467 ( .A(n12764), .B(n11985), .C(n14222), .Z(n14214) );
  HS65_LL_NAND2X2 U14468 ( .A(n11986), .B(n12103), .Z(n12768) );
  HS65_LL_NAND2X2 U14469 ( .A(n12768), .B(n14190), .Z(n14206) );
  HS65_LL_NAND4ABX3 U14470 ( .A(n14214), .B(n14206), .C(n12772), .D(n11987), 
        .Z(n13910) );
  HS65_LL_NOR3X1 U14471 ( .A(n11988), .B(n12778), .C(n13910), .Z(n11990) );
  HS65_LL_NAND2X2 U14472 ( .A(n12117), .B(n11989), .Z(n12754) );
  HS65_LL_NOR4ABX2 U14473 ( .A(n11990), .B(n14212), .C(n14211), .D(n12754), 
        .Z(n12135) );
  HS65_LL_NAND4ABX3 U14474 ( .A(n12750), .B(n12777), .C(n11991), .D(n12135), 
        .Z(n11994) );
  HS65_LL_AOI12X2 U14475 ( .A(n12119), .B(n12120), .C(n12108), .Z(n14874) );
  HS65_LL_NOR4ABX2 U14476 ( .A(n14874), .B(n11993), .C(n13905), .D(n11992), 
        .Z(n13918) );
  HS65_LL_NAND4ABX3 U14477 ( .A(n12113), .B(n11994), .C(n13918), .D(n12115), 
        .Z(n12001) );
  HS65_LL_NOR3X1 U14478 ( .A(n13164), .B(n12134), .C(n14209), .Z(n13145) );
  HS65_LL_OAI112X1 U14479 ( .A(n11996), .B(n12781), .C(n12762), .D(n11995), 
        .Z(n11997) );
  HS65_LL_NOR3X1 U14480 ( .A(n11998), .B(n13921), .C(n11997), .Z(n11999) );
  HS65_LL_NAND4ABX3 U14481 ( .A(n12786), .B(n14213), .C(n13145), .D(n11999), 
        .Z(n12000) );
  HS65_LL_MX41X4 U14482 ( .D0(n12003), .S0(n14899), .D1(n12002), .S1(n14891), 
        .D2(n12001), .S2(n14233), .D3(n12000), .S3(n14893), .Z(n15664) );
  HS65_LL_MUXI21X2 U14483 ( .D0(n15726), .D1(n15677), .S0(n15664), .Z(n15684)
         );
  HS65_LL_NAND2X2 U14484 ( .A(n12697), .B(n13106), .Z(n14580) );
  HS65_LL_NAND4ABX3 U14485 ( .A(n12702), .B(n12004), .C(n13096), .D(n14580), 
        .Z(n14604) );
  HS65_LL_NAND2X2 U14486 ( .A(n13106), .B(n12712), .Z(n12005) );
  HS65_LL_NAND4ABX3 U14487 ( .A(n12703), .B(n12731), .C(n12741), .D(n12005), 
        .Z(n14610) );
  HS65_LL_NAND3X2 U14488 ( .A(n13781), .B(n14592), .C(n15200), .Z(n13794) );
  HS65_LL_IVX2 U14489 ( .A(n13794), .Z(n15213) );
  HS65_LL_NOR2X2 U14490 ( .A(sa03[1]), .B(n12006), .Z(n12008) );
  HS65_LL_IVX2 U14491 ( .A(n14577), .Z(n12740) );
  HS65_LL_AOI12X2 U14492 ( .A(n14595), .B(n12007), .C(n14594), .Z(n13110) );
  HS65_LL_AOI112X2 U14493 ( .A(n12009), .B(n12008), .C(n12740), .D(n13110), 
        .Z(n12011) );
  HS65_LL_NOR4ABX2 U14494 ( .A(n12011), .B(n15217), .C(n13784), .D(n12010), 
        .Z(n12012) );
  HS65_LL_NAND4ABX3 U14495 ( .A(n13127), .B(n14610), .C(n15213), .D(n12012), 
        .Z(n12049) );
  HS65_LL_IVX2 U14496 ( .A(n15215), .Z(n12708) );
  HS65_LL_NAND3X2 U14497 ( .A(n15217), .B(n12708), .C(n14918), .Z(n13128) );
  HS65_LL_NAND2X2 U14498 ( .A(n14592), .B(n15200), .Z(n12015) );
  HS65_LL_NOR2X2 U14499 ( .A(n13095), .B(n14908), .Z(n12727) );
  HS65_LL_NOR3X1 U14500 ( .A(n14573), .B(n12028), .C(n12013), .Z(n12014) );
  HS65_LL_NAND4ABX3 U14501 ( .A(n13128), .B(n12015), .C(n12727), .D(n12014), 
        .Z(n12016) );
  HS65_LL_NOR3X1 U14502 ( .A(n12731), .B(n12017), .C(n12016), .Z(n14929) );
  HS65_LL_NOR2X2 U14503 ( .A(n12018), .B(n12711), .Z(n12725) );
  HS65_LL_OAI21X2 U14504 ( .A(n14594), .B(n14595), .C(n13772), .Z(n13783) );
  HS65_LL_NOR4ABX2 U14505 ( .A(n14929), .B(n12725), .C(n14917), .D(n13783), 
        .Z(n13768) );
  HS65_LL_IVX2 U14506 ( .A(n13773), .Z(n13779) );
  HS65_LL_NOR2X2 U14507 ( .A(n14595), .B(n13790), .Z(n12719) );
  HS65_LL_NOR2X2 U14508 ( .A(n12715), .B(n12719), .Z(n13775) );
  HS65_LL_NAND4ABX3 U14509 ( .A(n13779), .B(n14604), .C(n12019), .D(n13775), 
        .Z(n12020) );
  HS65_LL_NOR4ABX2 U14510 ( .A(n15214), .B(n13768), .C(n12021), .D(n12020), 
        .Z(n12047) );
  HS65_LL_IVX2 U14511 ( .A(n15240), .Z(n12046) );
  HS65_LL_NOR2X2 U14512 ( .A(n12022), .B(n14594), .Z(n12023) );
  HS65_LL_IVX2 U14513 ( .A(n15227), .Z(n12717) );
  HS65_LL_NAND4ABX3 U14514 ( .A(n12703), .B(n12023), .C(n12717), .D(n12036), 
        .Z(n14907) );
  HS65_LL_IVX2 U14515 ( .A(n15205), .Z(n12024) );
  HS65_LL_NAND2X2 U14516 ( .A(n14581), .B(n12024), .Z(n14596) );
  HS65_LL_OAI21X2 U14517 ( .A(n12026), .B(n12025), .C(n14571), .Z(n14606) );
  HS65_LL_AOI12X2 U14518 ( .A(n13790), .B(n12027), .C(n14925), .Z(n14566) );
  HS65_LL_NOR3X1 U14519 ( .A(n14596), .B(n14606), .C(n14566), .Z(n13770) );
  HS65_LL_AOI12X2 U14520 ( .A(n12712), .B(n13115), .C(n13094), .Z(n12032) );
  HS65_LL_NOR2AX3 U14521 ( .A(n15196), .B(n12028), .Z(n12734) );
  HS65_LL_NOR2X2 U14522 ( .A(n13113), .B(n14593), .Z(n14914) );
  HS65_LL_NAND3X2 U14523 ( .A(n12032), .B(n12734), .C(n14914), .Z(n12029) );
  HS65_LL_NOR4ABX2 U14524 ( .A(n13770), .B(n12741), .C(n14611), .D(n12029), 
        .Z(n15218) );
  HS65_LL_NAND4ABX3 U14525 ( .A(n13129), .B(n12030), .C(n15218), .D(n15200), 
        .Z(n12031) );
  HS65_LL_OAI13X1 U14526 ( .A(n14907), .B(n13110), .C(n12031), .D(n15234), .Z(
        n12045) );
  HS65_LL_OAI21X2 U14527 ( .A(n12696), .B(n13115), .C(n12697), .Z(n13100) );
  HS65_LL_NOR2X2 U14528 ( .A(n14595), .B(n13111), .Z(n14922) );
  HS65_LL_NOR2X2 U14529 ( .A(n12731), .B(n13108), .Z(n14565) );
  HS65_LL_NAND4ABX3 U14530 ( .A(n14921), .B(n12033), .C(n14565), .D(n12032), 
        .Z(n13124) );
  HS65_LL_NOR3X1 U14531 ( .A(n14922), .B(n14908), .C(n13124), .Z(n12034) );
  HS65_LL_IVX2 U14532 ( .A(n13129), .Z(n13786) );
  HS65_LL_NAND3X2 U14533 ( .A(n13100), .B(n12034), .C(n13786), .Z(n15226) );
  HS65_LL_NAND2X2 U14534 ( .A(n12035), .B(n12741), .Z(n12042) );
  HS65_LL_IVX2 U14535 ( .A(n12036), .Z(n14920) );
  HS65_LL_NOR2X2 U14536 ( .A(n14920), .B(n14573), .Z(n13116) );
  HS65_LL_NAND4ABX3 U14537 ( .A(n13774), .B(n13113), .C(n12730), .D(n13116), 
        .Z(n12041) );
  HS65_LL_OAI112X1 U14538 ( .A(n13790), .B(n12038), .C(n12037), .D(n13772), 
        .Z(n12039) );
  HS65_LL_NOR3X1 U14539 ( .A(n12715), .B(n13128), .C(n12039), .Z(n14587) );
  HS65_LL_NAND4ABX3 U14540 ( .A(n12042), .B(n12041), .C(n12040), .D(n14587), 
        .Z(n12043) );
  HS65_LL_OAI13X1 U14541 ( .A(n15226), .B(n14604), .C(n12043), .D(n15236), .Z(
        n12044) );
  HS65_LL_OAI112X1 U14542 ( .A(n12047), .B(n12046), .C(n12045), .D(n12044), 
        .Z(n12048) );
  HS65_LL_CBI4I6X2 U14543 ( .A(n14604), .B(n12049), .C(n15238), .D(n12048), 
        .Z(n15243) );
  HS65_LL_NOR2X2 U14544 ( .A(n12050), .B(n14707), .Z(n13720) );
  HS65_LL_NOR2X2 U14545 ( .A(n14723), .B(n13188), .Z(n12052) );
  HS65_LL_NAND2X2 U14546 ( .A(n12051), .B(n13722), .Z(n12081) );
  HS65_LL_NOR4ABX2 U14547 ( .A(n13720), .B(n12053), .C(n12052), .D(n12081), 
        .Z(n12099) );
  HS65_LL_NOR2X2 U14548 ( .A(n12055), .B(n12054), .Z(n12060) );
  HS65_LL_AOI13X2 U14549 ( .A(sa32[3]), .B(sa32[5]), .C(n12086), .D(n13287), 
        .Z(n12058) );
  HS65_LL_NAND2X2 U14550 ( .A(n12056), .B(n12086), .Z(n12057) );
  HS65_LL_NAND2X2 U14551 ( .A(n14357), .B(n14710), .Z(n14718) );
  HS65_LL_NAND4ABX3 U14552 ( .A(n14718), .B(n14706), .C(n14729), .D(n14728), 
        .Z(n13761) );
  HS65_LL_NOR4ABX2 U14553 ( .A(n12058), .B(n12057), .C(n13269), .D(n13761), 
        .Z(n12059) );
  HS65_LL_NAND3X2 U14554 ( .A(n12059), .B(n14364), .C(n12082), .Z(n14358) );
  HS65_LL_NOR4ABX2 U14555 ( .A(n12061), .B(n13279), .C(n12060), .D(n14358), 
        .Z(n12098) );
  HS65_LL_NAND2X2 U14556 ( .A(n13256), .B(n13277), .Z(n13738) );
  HS65_LL_NAND2X2 U14557 ( .A(n13266), .B(n13738), .Z(n13736) );
  HS65_LL_NAND2AX4 U14558 ( .A(n12062), .B(n14720), .Z(n13185) );
  HS65_LL_NOR4ABX2 U14559 ( .A(n13186), .B(n13193), .C(n12064), .D(n12063), 
        .Z(n14382) );
  HS65_LL_NAND2X2 U14560 ( .A(n14360), .B(n13178), .Z(n14699) );
  HS65_LL_NOR3AX2 U14561 ( .A(n12070), .B(n12065), .C(n14699), .Z(n12066) );
  HS65_LL_NAND4ABX3 U14562 ( .A(n13736), .B(n13185), .C(n14382), .D(n12066), 
        .Z(n12096) );
  HS65_LL_NOR4ABX2 U14563 ( .A(n14737), .B(n12077), .C(n13256), .D(n12083), 
        .Z(n12069) );
  HS65_LL_NAND3X2 U14564 ( .A(n14720), .B(n12067), .C(n14361), .Z(n14370) );
  HS65_LL_NOR4ABX2 U14565 ( .A(n12070), .B(n12069), .C(n12068), .D(n14370), 
        .Z(n12094) );
  HS65_LL_NOR2X2 U14566 ( .A(n13258), .B(n12071), .Z(n12072) );
  HS65_LL_NAND4ABX3 U14567 ( .A(n13181), .B(n12073), .C(n12072), .D(n13264), 
        .Z(n12092) );
  HS65_LL_AOI12X2 U14568 ( .A(n12086), .B(n14733), .C(n12074), .Z(n13184) );
  HS65_LL_NOR4ABX2 U14569 ( .A(n13184), .B(n12076), .C(n13257), .D(n12075), 
        .Z(n12078) );
  HS65_LL_NAND4ABX3 U14570 ( .A(n13275), .B(n12079), .C(n12078), .D(n12077), 
        .Z(n14717) );
  HS65_LL_IVX2 U14571 ( .A(n12080), .Z(n13249) );
  HS65_LL_NAND3X2 U14572 ( .A(n13718), .B(n14372), .C(n13249), .Z(n14359) );
  HS65_LL_NOR3X1 U14573 ( .A(n14735), .B(n14359), .C(n12081), .Z(n13747) );
  HS65_LL_NAND4ABX3 U14574 ( .A(n12084), .B(n12083), .C(n13747), .D(n12082), 
        .Z(n12085) );
  HS65_LL_AOI12X2 U14575 ( .A(n12087), .B(n12086), .C(n12085), .Z(n13260) );
  HS65_LL_NAND4ABX3 U14576 ( .A(n12089), .B(n14717), .C(n13260), .D(n12088), 
        .Z(n12090) );
  HS65_LL_OAI13X1 U14577 ( .A(n12092), .B(n12091), .C(n12090), .D(n14742), .Z(
        n12093) );
  HS65_LL_CBI4I1X3 U14578 ( .A(n13746), .B(n12094), .C(n13744), .D(n12093), 
        .Z(n12095) );
  HS65_LL_CBI4I6X2 U14579 ( .A(n14727), .B(n12096), .C(n14748), .D(n12095), 
        .Z(n12097) );
  HS65_LL_CBI4I1X3 U14580 ( .A(n12099), .B(n12098), .C(n14380), .D(n12097), 
        .Z(n15701) );
  HS65_LL_MUXI21X2 U14581 ( .D0(n15242), .D1(w3[29]), .S0(n15701), .Z(n12100)
         );
  HS65_LLS_XOR3X2 U14582 ( .A(n15684), .B(n15243), .C(n12100), .Z(n12147) );
  HS65_LL_NAND3AX3 U14583 ( .A(n12101), .B(n12111), .C(n12768), .Z(n14200) );
  HS65_LL_IVX2 U14584 ( .A(n12799), .Z(n14208) );
  HS65_LL_NAND3X2 U14585 ( .A(n12770), .B(n14208), .C(n14886), .Z(n12133) );
  HS65_LL_NOR2X2 U14586 ( .A(n12777), .B(n12102), .Z(n13152) );
  HS65_LL_NAND2X2 U14587 ( .A(n12103), .B(n14196), .Z(n14867) );
  HS65_LL_NAND3X2 U14588 ( .A(n13152), .B(n12104), .C(n14867), .Z(n14189) );
  HS65_LL_NAND4ABX3 U14589 ( .A(n13163), .B(n12780), .C(n12105), .D(n14188), 
        .Z(n12106) );
  HS65_LL_NOR4ABX2 U14590 ( .A(n13145), .B(n12794), .C(n14189), .D(n12106), 
        .Z(n12107) );
  HS65_LL_NAND4ABX3 U14591 ( .A(n12108), .B(n12133), .C(n12107), .D(n13915), 
        .Z(n12143) );
  HS65_LL_IVX2 U14592 ( .A(n12109), .Z(n13922) );
  HS65_LL_NOR4ABX2 U14593 ( .A(n12111), .B(n12110), .C(n13922), .D(n14189), 
        .Z(n12141) );
  HS65_LL_NOR2X2 U14594 ( .A(n14221), .B(n12112), .Z(n13165) );
  HS65_LL_NOR2X2 U14595 ( .A(n12114), .B(n12113), .Z(n13144) );
  HS65_LL_IVX2 U14596 ( .A(n13144), .Z(n12125) );
  HS65_LL_NAND2X2 U14597 ( .A(n12761), .B(n13913), .Z(n13925) );
  HS65_LL_NOR4ABX2 U14598 ( .A(n12116), .B(n12115), .C(n12125), .D(n13925), 
        .Z(n14226) );
  HS65_LL_NAND2X2 U14599 ( .A(n14226), .B(n12803), .Z(n13161) );
  HS65_LL_NAND2AX4 U14600 ( .A(n14219), .B(n12117), .Z(n14878) );
  HS65_LL_NOR4ABX2 U14601 ( .A(n13165), .B(n12118), .C(n13161), .D(n14878), 
        .Z(n12140) );
  HS65_LL_AOI12X2 U14602 ( .A(n12120), .B(n12119), .C(n12787), .Z(n13930) );
  HS65_LL_NAND2X2 U14603 ( .A(n13924), .B(n13923), .Z(n12124) );
  HS65_LL_NOR4ABX2 U14604 ( .A(n12122), .B(n14220), .C(n14221), .D(n12121), 
        .Z(n12123) );
  HS65_LL_NAND4ABX3 U14605 ( .A(n12125), .B(n12124), .C(n13145), .D(n12123), 
        .Z(n14875) );
  HS65_LL_NAND4ABX3 U14606 ( .A(n12799), .B(n12780), .C(n12760), .D(n13913), 
        .Z(n12126) );
  HS65_LL_NOR3X1 U14607 ( .A(n13148), .B(n14875), .C(n12126), .Z(n13907) );
  HS65_LL_NAND4ABX3 U14608 ( .A(n12127), .B(n13156), .C(n13930), .D(n13907), 
        .Z(n12130) );
  HS65_LL_NAND4ABX3 U14609 ( .A(n14189), .B(n12130), .C(n12129), .D(n12128), 
        .Z(n12138) );
  HS65_LL_NAND2X2 U14610 ( .A(n12131), .B(n13923), .Z(n12797) );
  HS65_LL_AOI12X2 U14611 ( .A(n12132), .B(n12788), .C(n12797), .Z(n14865) );
  HS65_LL_NOR4ABX2 U14612 ( .A(n12135), .B(n13916), .C(n12134), .D(n12133), 
        .Z(n12136) );
  HS65_LL_AOI13X2 U14613 ( .A(n14865), .B(n14203), .C(n12136), .D(n12774), .Z(
        n12137) );
  HS65_LL_CBI4I6X2 U14614 ( .A(n14213), .B(n12138), .C(n14891), .D(n12137), 
        .Z(n12139) );
  HS65_LL_CBI4I1X3 U14615 ( .A(n12141), .B(n12140), .C(n14895), .D(n12139), 
        .Z(n12142) );
  HS65_LL_CBI4I6X2 U14616 ( .A(n14200), .B(n12143), .C(n14893), .D(n12142), 
        .Z(n15338) );
  HS65_LL_OAI21X2 U14617 ( .A(n15338), .B(n12147), .C(n14808), .Z(n12146) );
  HS65_LL_IVX2 U14618 ( .A(text_in_r[29]), .Z(n12144) );
  HS65_LL_OAI212X3 U14619 ( .A(w3[29]), .B(text_in_r[29]), .C(n15242), .D(
        n12144), .E(n15545), .Z(n12145) );
  HS65_LL_CBI4I1X3 U14620 ( .A(n12147), .B(n15338), .C(n12146), .D(n12145), 
        .Z(N87) );
  HS65_LLS_XNOR2X3 U14621 ( .A(n12148), .B(n15127), .Z(n14984) );
  HS65_LL_OAI112X1 U14622 ( .A(n12151), .B(n12150), .C(n12149), .D(n12827), 
        .Z(n12152) );
  HS65_LL_NOR4ABX2 U14623 ( .A(n12154), .B(n12811), .C(n12153), .D(n12152), 
        .Z(n12155) );
  HS65_LL_NAND4ABX3 U14624 ( .A(n12820), .B(n14669), .C(n12175), .D(n12155), 
        .Z(n12193) );
  HS65_LL_NOR4ABX2 U14625 ( .A(n12158), .B(n12157), .C(n14661), .D(n12156), 
        .Z(n12159) );
  HS65_LL_NAND4ABX3 U14626 ( .A(n12181), .B(n12160), .C(n12816), .D(n12159), 
        .Z(n12191) );
  HS65_LL_NAND3X2 U14627 ( .A(n12162), .B(n12830), .C(n12161), .Z(n14668) );
  HS65_LL_NAND4ABX3 U14628 ( .A(n14661), .B(n14668), .C(n12164), .D(n12163), 
        .Z(n12171) );
  HS65_LL_CBI4I6X2 U14629 ( .A(n12168), .B(n12167), .C(n12166), .D(n12165), 
        .Z(n12170) );
  HS65_LL_NOR4ABX2 U14630 ( .A(n12170), .B(n12169), .C(n14657), .D(n12826), 
        .Z(n14677) );
  HS65_LL_NAND4ABX3 U14631 ( .A(n12819), .B(n12171), .C(n12175), .D(n14677), 
        .Z(n12190) );
  HS65_LL_NAND2X2 U14632 ( .A(n12173), .B(n12172), .Z(n14656) );
  HS65_LL_NAND3X2 U14633 ( .A(n12175), .B(n12174), .C(n12829), .Z(n12188) );
  HS65_LL_NOR2X2 U14634 ( .A(n12846), .B(n12176), .Z(n12187) );
  HS65_LL_NAND2X2 U14635 ( .A(n12178), .B(n12177), .Z(n12179) );
  HS65_LL_NOR3X1 U14636 ( .A(n12181), .B(n12180), .C(n12179), .Z(n12185) );
  HS65_LL_NOR4ABX2 U14637 ( .A(n12185), .B(n12184), .C(n12183), .D(n12182), 
        .Z(n12186) );
  HS65_LL_NAND4ABX3 U14638 ( .A(n14656), .B(n12188), .C(n12187), .D(n12186), 
        .Z(n12189) );
  HS65_LL_MX41X4 U14639 ( .D0(n12193), .S0(n12192), .D1(n12191), .S1(n14691), 
        .D2(n12190), .S2(n14683), .D3(n12189), .S3(n14685), .Z(n14837) );
  HS65_LL_IVX2 U14640 ( .A(n14837), .Z(n15447) );
  HS65_LL_MUXI21X2 U14641 ( .D0(n14837), .D1(n15447), .S0(w1[13]), .Z(n12194)
         );
  HS65_LLS_XOR3X2 U14642 ( .A(n14984), .B(n12194), .C(n15267), .Z(n12236) );
  HS65_LL_NOR3AX2 U14643 ( .A(n12196), .B(n13429), .C(n12195), .Z(n12198) );
  HS65_LL_NAND3X2 U14644 ( .A(n12199), .B(n12198), .C(n12197), .Z(n13426) );
  HS65_LL_AOI12X2 U14645 ( .A(n12202), .B(n12201), .C(n12200), .Z(n13413) );
  HS65_LL_NAND2X2 U14646 ( .A(n12203), .B(n13417), .Z(n14298) );
  HS65_LL_NOR4ABX2 U14647 ( .A(n14323), .B(n13413), .C(n12226), .D(n14298), 
        .Z(n12204) );
  HS65_LL_NAND4ABX3 U14648 ( .A(n12205), .B(n14319), .C(n14330), .D(n12204), 
        .Z(n12232) );
  HS65_LL_NAND4ABX3 U14649 ( .A(n13433), .B(n12207), .C(n12206), .D(n14293), 
        .Z(n12208) );
  HS65_LL_NOR4ABX2 U14650 ( .A(n12216), .B(n12210), .C(n12209), .D(n12208), 
        .Z(n12230) );
  HS65_LL_NOR2X2 U14651 ( .A(n12212), .B(n12211), .Z(n12214) );
  HS65_LL_NOR4ABX2 U14652 ( .A(n14315), .B(n12214), .C(n12213), .D(n14292), 
        .Z(n12215) );
  HS65_LL_NAND4ABX3 U14653 ( .A(n12217), .B(n13432), .C(n12216), .D(n12215), 
        .Z(n12218) );
  HS65_LL_OAI13X1 U14654 ( .A(n12226), .B(n13456), .C(n12218), .D(n14339), .Z(
        n12228) );
  HS65_LL_NOR3X1 U14655 ( .A(n12220), .B(n14304), .C(n12219), .Z(n12221) );
  HS65_LL_NAND4ABX3 U14656 ( .A(n12223), .B(n13421), .C(n12222), .D(n12221), 
        .Z(n12224) );
  HS65_LL_OAI13X1 U14657 ( .A(n12226), .B(n12225), .C(n12224), .D(n14335), .Z(
        n12227) );
  HS65_LL_OAI112X1 U14658 ( .A(n12230), .B(n12229), .C(n12228), .D(n12227), 
        .Z(n12231) );
  HS65_LL_CBI4I6X2 U14659 ( .A(n13426), .B(n12232), .C(n14337), .D(n12231), 
        .Z(n15363) );
  HS65_LL_OAI21X2 U14660 ( .A(n15363), .B(n12236), .C(n14832), .Z(n12235) );
  HS65_LL_IVX2 U14661 ( .A(text_in_r[77]), .Z(n12233) );
  HS65_LL_OAI212X3 U14662 ( .A(w1[13]), .B(text_in_r[77]), .C(n15362), .D(
        n12233), .E(n15545), .Z(n12234) );
  HS65_LL_CBI4I1X3 U14663 ( .A(n12236), .B(n15363), .C(n12235), .D(n12234), 
        .Z(N183) );
  HS65_LL_IVX2 U14664 ( .A(n15425), .Z(n15426) );
  HS65_LL_MUXI21X2 U14665 ( .D0(n15425), .D1(n15426), .S0(w2[17]), .Z(n12346)
         );
  HS65_LL_NAND3X2 U14666 ( .A(n12237), .B(n15291), .C(n12260), .Z(n12246) );
  HS65_LL_NOR4ABX2 U14667 ( .A(n15311), .B(n12239), .C(n12278), .D(n12238), 
        .Z(n12241) );
  HS65_LL_NOR4ABX2 U14668 ( .A(n12242), .B(n12241), .C(n12240), .D(n14514), 
        .Z(n14524) );
  HS65_LL_NOR3X1 U14669 ( .A(n12244), .B(n14503), .C(n12243), .Z(n12245) );
  HS65_LL_NAND4ABX3 U14670 ( .A(n12247), .B(n12246), .C(n14524), .D(n12245), 
        .Z(n12292) );
  HS65_LL_NOR2X2 U14671 ( .A(n15303), .B(n12248), .Z(n12254) );
  HS65_LL_NOR3AX2 U14672 ( .A(n12250), .B(n12249), .C(n14514), .Z(n14529) );
  HS65_LL_NAND3X2 U14673 ( .A(n12269), .B(n12260), .C(n12251), .Z(n12252) );
  HS65_LL_NOR4ABX2 U14674 ( .A(n12254), .B(n14529), .C(n12253), .D(n12252), 
        .Z(n12255) );
  HS65_LL_NAND3X2 U14675 ( .A(n12256), .B(n15288), .C(n12255), .Z(n12291) );
  HS65_LL_NOR3X1 U14676 ( .A(n12258), .B(n14526), .C(n12257), .Z(n14508) );
  HS65_LL_IVX2 U14677 ( .A(n12259), .Z(n12261) );
  HS65_LL_NAND2X2 U14678 ( .A(n12261), .B(n12260), .Z(n15306) );
  HS65_LL_AOI112X2 U14679 ( .A(n12264), .B(n12263), .C(n12262), .D(n15306), 
        .Z(n12267) );
  HS65_LL_NOR4ABX2 U14680 ( .A(n12267), .B(n12266), .C(n12288), .D(n12265), 
        .Z(n12268) );
  HS65_LL_NAND3X2 U14681 ( .A(n12269), .B(n14508), .C(n12268), .Z(n12290) );
  HS65_LL_NAND2X2 U14682 ( .A(n12271), .B(n12270), .Z(n12282) );
  HS65_LL_OAI112X1 U14683 ( .A(sa13[7]), .B(n12274), .C(n12273), .D(n12272), 
        .Z(n12275) );
  HS65_LL_NOR4ABX2 U14684 ( .A(n12277), .B(n12276), .C(n15317), .D(n12275), 
        .Z(n15309) );
  HS65_LL_NOR4ABX2 U14685 ( .A(n12280), .B(n12279), .C(n12278), .D(n14515), 
        .Z(n12281) );
  HS65_LL_NAND4ABX3 U14686 ( .A(n12283), .B(n12282), .C(n15309), .D(n12281), 
        .Z(n12287) );
  HS65_LL_NOR2X2 U14687 ( .A(n12285), .B(n12284), .Z(n14532) );
  HS65_LL_NAND4ABX3 U14688 ( .A(n12288), .B(n12287), .C(n12286), .D(n14532), 
        .Z(n12289) );
  HS65_LL_MX41X4 U14689 ( .D0(n12292), .S0(n15328), .D1(n12291), .S1(n15326), 
        .D2(n12290), .S2(n15324), .D3(n12289), .S3(n15322), .Z(n15599) );
  HS65_LL_IVX2 U14690 ( .A(n15599), .Z(n15336) );
  HS65_LL_IVX2 U14691 ( .A(n12318), .Z(n12295) );
  HS65_LL_NAND4ABX3 U14692 ( .A(n15376), .B(n12295), .C(n12294), .D(n12293), 
        .Z(n12298) );
  HS65_LL_NAND4ABX3 U14693 ( .A(n12299), .B(n12298), .C(n12297), .D(n12296), 
        .Z(n12345) );
  HS65_LL_NOR4ABX2 U14694 ( .A(n12303), .B(n12302), .C(n12301), .D(n12300), 
        .Z(n12304) );
  HS65_LL_NAND4ABX3 U14695 ( .A(n12307), .B(n12306), .C(n12305), .D(n12304), 
        .Z(n15387) );
  HS65_LL_NOR2X2 U14696 ( .A(n12308), .B(n13040), .Z(n12312) );
  HS65_LL_NOR4ABX2 U14697 ( .A(n12312), .B(n12311), .C(n12310), .D(n12309), 
        .Z(n12320) );
  HS65_LL_NAND3AX3 U14698 ( .A(n12315), .B(n12314), .C(n12313), .Z(n13026) );
  HS65_LL_NOR4ABX2 U14699 ( .A(n12318), .B(n12317), .C(n12316), .D(n13026), 
        .Z(n12319) );
  HS65_LL_NAND4ABX3 U14700 ( .A(n12321), .B(n15387), .C(n12320), .D(n12319), 
        .Z(n12344) );
  HS65_LL_NAND4ABX3 U14701 ( .A(n12323), .B(n13034), .C(n13025), .D(n12322), 
        .Z(n12329) );
  HS65_LL_NOR4ABX2 U14702 ( .A(n12326), .B(n12325), .C(n12324), .D(n15376), 
        .Z(n12327) );
  HS65_LL_NAND4ABX3 U14703 ( .A(n15402), .B(n12329), .C(n12328), .D(n12327), 
        .Z(n12343) );
  HS65_LL_AND2X4 U14704 ( .A(n15392), .B(n15393), .Z(n12339) );
  HS65_LL_NOR4ABX2 U14705 ( .A(n12332), .B(n12331), .C(n13034), .D(n12330), 
        .Z(n12333) );
  HS65_LL_NAND3X2 U14706 ( .A(n12334), .B(n15391), .C(n12333), .Z(n13018) );
  HS65_LL_NOR4ABX2 U14707 ( .A(n12337), .B(n12336), .C(n12335), .D(n13018), 
        .Z(n12338) );
  HS65_LL_NAND4ABX3 U14708 ( .A(n12341), .B(n12340), .C(n12339), .D(n12338), 
        .Z(n12342) );
  HS65_LL_MX41X4 U14709 ( .D0(n12345), .S0(n13020), .D1(n12344), .S1(n15416), 
        .D2(n12343), .S2(n15408), .D3(n12342), .S3(n15400), .Z(n15578) );
  HS65_LL_MUXI21X2 U14710 ( .D0(n15599), .D1(n15336), .S0(n15578), .Z(n15623)
         );
  HS65_LLS_XOR3X2 U14711 ( .A(n15579), .B(n12346), .C(n15623), .Z(n12392) );
  HS65_LL_NOR4ABX2 U14712 ( .A(n12349), .B(n12348), .C(n13335), .D(n12347), 
        .Z(n13078) );
  HS65_LL_NOR2AX3 U14713 ( .A(n12351), .B(n12350), .Z(n15490) );
  HS65_LL_NAND2X2 U14714 ( .A(n12352), .B(n15482), .Z(n13054) );
  HS65_LL_NOR4ABX2 U14715 ( .A(n15490), .B(n12353), .C(n12384), .D(n13054), 
        .Z(n12354) );
  HS65_LL_NAND3X2 U14716 ( .A(n13078), .B(n12355), .C(n12354), .Z(n12388) );
  HS65_LL_NAND3X2 U14717 ( .A(n12358), .B(n12357), .C(n12356), .Z(n13069) );
  HS65_LL_AOI112X2 U14718 ( .A(sa31[7]), .B(n12360), .C(sa31[6]), .D(n12359), 
        .Z(n12361) );
  HS65_LL_NOR4ABX2 U14719 ( .A(n12363), .B(n13344), .C(n12362), .D(n12361), 
        .Z(n12364) );
  HS65_LL_NAND4ABX3 U14720 ( .A(n13079), .B(n13069), .C(n13334), .D(n12364), 
        .Z(n12387) );
  HS65_LL_NOR2X2 U14721 ( .A(n12377), .B(n13310), .Z(n13342) );
  HS65_LL_NAND4ABX3 U14722 ( .A(n12366), .B(n15481), .C(n12365), .D(n13342), 
        .Z(n12368) );
  HS65_LL_NAND4ABX3 U14723 ( .A(n15505), .B(n12368), .C(n13327), .D(n12367), 
        .Z(n12386) );
  HS65_LL_NOR3X1 U14724 ( .A(sa31[7]), .B(n12370), .C(n12369), .Z(n15477) );
  HS65_LL_NAND3AX3 U14725 ( .A(n12372), .B(n12371), .C(n13325), .Z(n12373) );
  HS65_LL_NOR3X1 U14726 ( .A(n12374), .B(n15477), .C(n12373), .Z(n13071) );
  HS65_LL_NOR2X2 U14727 ( .A(n12376), .B(n12375), .Z(n13055) );
  HS65_LL_NOR3X1 U14728 ( .A(n12378), .B(n12377), .C(n13055), .Z(n15474) );
  HS65_LL_NAND2X2 U14729 ( .A(n12379), .B(n13347), .Z(n13075) );
  HS65_LL_NOR4ABX2 U14730 ( .A(n15474), .B(n12381), .C(n12380), .D(n13075), 
        .Z(n12382) );
  HS65_LL_NAND4ABX3 U14731 ( .A(n12384), .B(n12383), .C(n13071), .D(n12382), 
        .Z(n12385) );
  HS65_LL_MX41X4 U14732 ( .D0(n12388), .S0(n15478), .D1(n12387), .S1(n15494), 
        .D2(n12386), .S2(n13352), .D3(n12385), .S3(n15503), .Z(n15511) );
  HS65_LLS_XOR2X3 U14733 ( .A(n15511), .B(n15192), .Z(n15631) );
  HS65_LL_OAI21X2 U14734 ( .A(n15631), .B(n12392), .C(n14832), .Z(n12391) );
  HS65_LL_AOI12X2 U14735 ( .A(w2[17]), .B(text_in_r[49]), .C(n14808), .Z(
        n12389) );
  HS65_LL_OAI21X2 U14736 ( .A(w2[17]), .B(text_in_r[49]), .C(n12389), .Z(
        n12390) );
  HS65_LL_CBI4I1X3 U14737 ( .A(n12392), .B(n15631), .C(n12391), .D(n12390), 
        .Z(N131) );
  HS65_LL_NAND4ABX3 U14738 ( .A(n12395), .B(n13971), .C(n12394), .D(n12393), 
        .Z(n12396) );
  HS65_LL_NAND4ABX3 U14739 ( .A(n12997), .B(n12396), .C(n13581), .D(n13958), 
        .Z(n12437) );
  HS65_LL_NOR3X1 U14740 ( .A(n12398), .B(n13598), .C(n12397), .Z(n12991) );
  HS65_LL_NAND3X2 U14741 ( .A(n12400), .B(n12399), .C(n13953), .Z(n12402) );
  HS65_LL_NAND4ABX3 U14742 ( .A(n12978), .B(n12402), .C(n12401), .D(n13581), 
        .Z(n13947) );
  HS65_LL_NOR3X1 U14743 ( .A(n12413), .B(n12412), .C(n13947), .Z(n12404) );
  HS65_LL_NAND4ABX3 U14744 ( .A(n13576), .B(n12999), .C(n12404), .D(n12403), 
        .Z(n13567) );
  HS65_LL_NAND4ABX3 U14745 ( .A(n12407), .B(n13567), .C(n12406), .D(n12405), 
        .Z(n12408) );
  HS65_LL_NOR4ABX2 U14746 ( .A(n12411), .B(n12410), .C(n12409), .D(n12408), 
        .Z(n12435) );
  HS65_LL_NOR2X2 U14747 ( .A(n12413), .B(n12412), .Z(n12414) );
  HS65_LL_NAND4ABX3 U14748 ( .A(n12416), .B(n12415), .C(n12414), .D(n13593), 
        .Z(n12420) );
  HS65_LL_NOR2X2 U14749 ( .A(n13583), .B(n13574), .Z(n13944) );
  HS65_LL_NOR4ABX2 U14750 ( .A(n13944), .B(n12418), .C(n12962), .D(n12417), 
        .Z(n13000) );
  HS65_LL_NAND4ABX3 U14751 ( .A(n12421), .B(n12420), .C(n12419), .D(n13000), 
        .Z(n12432) );
  HS65_LL_NAND2X2 U14752 ( .A(n12423), .B(n12422), .Z(n13570) );
  HS65_LL_NOR3X1 U14753 ( .A(n13599), .B(n12424), .C(n13570), .Z(n12426) );
  HS65_LL_NOR4ABX2 U14754 ( .A(n12427), .B(n12426), .C(n12425), .D(n12969), 
        .Z(n12428) );
  HS65_LL_NAND3X2 U14755 ( .A(n12430), .B(n12429), .C(n12428), .Z(n12431) );
  HS65_LL_AOI22X1 U14756 ( .A(n13981), .B(n12432), .C(n13972), .D(n12431), .Z(
        n12433) );
  HS65_LL_CBI4I1X3 U14757 ( .A(n12991), .B(n12435), .C(n12434), .D(n12433), 
        .Z(n12436) );
  HS65_LL_CBI4I6X2 U14758 ( .A(n13955), .B(n12437), .C(n13614), .D(n12436), 
        .Z(n15256) );
  HS65_LL_NAND4ABX3 U14759 ( .A(n12439), .B(n12438), .C(n12533), .D(n12447), 
        .Z(n12445) );
  HS65_LL_NOR4ABX2 U14760 ( .A(n12443), .B(n12442), .C(n12441), .D(n12440), 
        .Z(n12444) );
  HS65_LL_NAND4ABX3 U14761 ( .A(n12513), .B(n12445), .C(n12949), .D(n12444), 
        .Z(n12484) );
  HS65_LL_NOR2X2 U14762 ( .A(n12446), .B(n12928), .Z(n12491) );
  HS65_LL_NAND2X2 U14763 ( .A(n12448), .B(n12447), .Z(n12912) );
  HS65_LL_NAND4ABX3 U14764 ( .A(n12451), .B(n12912), .C(n12450), .D(n12449), 
        .Z(n12452) );
  HS65_LL_NOR4ABX2 U14765 ( .A(n12454), .B(n12491), .C(n12453), .D(n12452), 
        .Z(n12455) );
  HS65_LL_NAND3X2 U14766 ( .A(n12457), .B(n12456), .C(n12455), .Z(n12483) );
  HS65_LL_IVX2 U14767 ( .A(n12458), .Z(n12493) );
  HS65_LL_NAND4ABX3 U14768 ( .A(n12460), .B(n12493), .C(n12459), .D(n12533), 
        .Z(n12940) );
  HS65_LL_NAND4ABX3 U14769 ( .A(n12462), .B(n12492), .C(n12470), .D(n12461), 
        .Z(n12465) );
  HS65_LL_NAND4ABX3 U14770 ( .A(n12940), .B(n12465), .C(n12464), .D(n12463), 
        .Z(n12482) );
  HS65_LL_NAND4ABX3 U14771 ( .A(n12469), .B(n12468), .C(n12467), .D(n12466), 
        .Z(n12497) );
  HS65_LL_IVX2 U14772 ( .A(n12470), .Z(n12486) );
  HS65_LL_NOR3X1 U14773 ( .A(n12486), .B(n12472), .C(n12471), .Z(n12474) );
  HS65_LL_NAND3X2 U14774 ( .A(n12475), .B(n12474), .C(n12473), .Z(n12525) );
  HS65_LL_NOR4ABX2 U14775 ( .A(n12478), .B(n12477), .C(n12476), .D(n12525), 
        .Z(n12479) );
  HS65_LL_NAND4ABX3 U14776 ( .A(n12913), .B(n12497), .C(n12480), .D(n12479), 
        .Z(n12481) );
  HS65_LL_MX41X4 U14777 ( .D0(n12484), .S0(n12540), .D1(n12483), .S1(n12951), 
        .D2(n12482), .S2(n12943), .D3(n12481), .S3(n12945), .Z(n15351) );
  HS65_LLS_XNOR2X3 U14778 ( .A(n15256), .B(n15351), .Z(n14831) );
  HS65_LL_NOR2X2 U14779 ( .A(n12486), .B(n12485), .Z(n12507) );
  HS65_LL_NOR4ABX2 U14780 ( .A(n12507), .B(n12489), .C(n12488), .D(n12487), 
        .Z(n12490) );
  HS65_LL_NAND4ABX3 U14781 ( .A(n12493), .B(n12492), .C(n12491), .D(n12490), 
        .Z(n12496) );
  HS65_LL_NAND4ABX3 U14782 ( .A(n12529), .B(n12496), .C(n12495), .D(n12494), 
        .Z(n12541) );
  HS65_LL_AOI112X2 U14783 ( .A(n12500), .B(n12499), .C(n12498), .D(n12497), 
        .Z(n12502) );
  HS65_LL_NAND4ABX3 U14784 ( .A(n12504), .B(n12503), .C(n12502), .D(n12501), 
        .Z(n12941) );
  HS65_LL_NOR4ABX2 U14785 ( .A(n12507), .B(n12506), .C(n12505), .D(n12941), 
        .Z(n12508) );
  HS65_LL_NAND4ABX3 U14786 ( .A(n12511), .B(n12510), .C(n12509), .D(n12508), 
        .Z(n12539) );
  HS65_LL_NOR3X1 U14787 ( .A(n12514), .B(n12513), .C(n12512), .Z(n12520) );
  HS65_LL_NOR4ABX2 U14788 ( .A(n12527), .B(n12515), .C(n12526), .D(n12937), 
        .Z(n12517) );
  HS65_LL_NAND3X2 U14789 ( .A(n12518), .B(n12517), .C(n12516), .Z(n12953) );
  HS65_LL_NOR4ABX2 U14790 ( .A(n12521), .B(n12520), .C(n12519), .D(n12953), 
        .Z(n12523) );
  HS65_LL_IVX2 U14791 ( .A(n12530), .Z(n12522) );
  HS65_LL_NAND4ABX3 U14792 ( .A(n12524), .B(n12529), .C(n12523), .D(n12522), 
        .Z(n12538) );
  HS65_LL_NOR4ABX2 U14793 ( .A(n12528), .B(n12527), .C(n12526), .D(n12525), 
        .Z(n12532) );
  HS65_LL_NOR4ABX2 U14794 ( .A(n12532), .B(n12531), .C(n12530), .D(n12529), 
        .Z(n12534) );
  HS65_LL_NAND4ABX3 U14795 ( .A(n12536), .B(n12535), .C(n12534), .D(n12533), 
        .Z(n12537) );
  HS65_LL_MX41X4 U14796 ( .D0(n12541), .S0(n12540), .D1(n12539), .S1(n12951), 
        .D2(n12538), .S2(n12943), .D3(n12537), .S3(n12945), .Z(n15543) );
  HS65_LL_MUXI21X2 U14797 ( .D0(w0[20]), .D1(n15255), .S0(n15543), .Z(n12542)
         );
  HS65_LLS_XOR3X2 U14798 ( .A(n14831), .B(n12542), .C(n13855), .Z(n12641) );
  HS65_LL_NAND2AX4 U14799 ( .A(n14002), .B(n12543), .Z(n13691) );
  HS65_LL_NAND2X2 U14800 ( .A(n12545), .B(n12544), .Z(n12567) );
  HS65_LL_NOR2X2 U14801 ( .A(n14000), .B(n12567), .Z(n13491) );
  HS65_LL_NOR3X1 U14802 ( .A(n13697), .B(n12546), .C(n14025), .Z(n14117) );
  HS65_LL_IVX2 U14803 ( .A(n13662), .Z(n12547) );
  HS65_LL_NOR2X2 U14804 ( .A(n12548), .B(n12547), .Z(n12551) );
  HS65_LL_NOR4ABX2 U14805 ( .A(n12551), .B(n12550), .C(n12584), .D(n12549), 
        .Z(n12888) );
  HS65_LL_NOR4ABX2 U14806 ( .A(n14117), .B(n12888), .C(n14004), .D(n13478), 
        .Z(n12552) );
  HS65_LL_NAND4ABX3 U14807 ( .A(n12553), .B(n13691), .C(n13491), .D(n12552), 
        .Z(n12595) );
  HS65_LL_NAND3AX3 U14808 ( .A(n14000), .B(n14114), .C(n12871), .Z(n14110) );
  HS65_LL_NOR2X2 U14809 ( .A(n12555), .B(n12554), .Z(n12556) );
  HS65_LL_NOR3X1 U14810 ( .A(n13687), .B(n12556), .C(n12891), .Z(n12566) );
  HS65_LL_NOR2X2 U14811 ( .A(n14094), .B(n13497), .Z(n12569) );
  HS65_LL_NAND2X2 U14812 ( .A(n13685), .B(n13662), .Z(n14011) );
  HS65_LL_NAND3AX3 U14813 ( .A(n14104), .B(n13489), .C(n12894), .Z(n13700) );
  HS65_LL_NAND3AX3 U14814 ( .A(n13700), .B(n12558), .C(n12557), .Z(n12559) );
  HS65_LL_NOR4ABX2 U14815 ( .A(n12560), .B(n12569), .C(n14011), .D(n12559), 
        .Z(n13993) );
  HS65_LL_NOR3X1 U14816 ( .A(n12562), .B(n14105), .C(n12561), .Z(n12563) );
  HS65_LL_NAND3X2 U14817 ( .A(n13670), .B(n13993), .C(n12563), .Z(n13675) );
  HS65_LL_NOR4ABX2 U14818 ( .A(n14103), .B(n13996), .C(n12564), .D(n13675), 
        .Z(n12565) );
  HS65_LL_NAND4ABX3 U14819 ( .A(n14110), .B(n12567), .C(n12566), .D(n12565), 
        .Z(n12594) );
  HS65_LL_NAND2AX4 U14820 ( .A(n14025), .B(n14111), .Z(n12571) );
  HS65_LL_NAND4ABX3 U14821 ( .A(n14105), .B(n13700), .C(n13491), .D(n13488), 
        .Z(n12570) );
  HS65_LL_NOR2AX3 U14822 ( .A(n13685), .B(n12568), .Z(n13498) );
  HS65_LL_NAND4ABX3 U14823 ( .A(n12571), .B(n12570), .C(n13498), .D(n12569), 
        .Z(n12575) );
  HS65_LL_NOR2X2 U14824 ( .A(n14096), .B(n13467), .Z(n12574) );
  HS65_LL_NOR2X2 U14825 ( .A(n14108), .B(n12572), .Z(n12573) );
  HS65_LL_NOR3X1 U14826 ( .A(n13672), .B(n12874), .C(n12573), .Z(n13475) );
  HS65_LL_NAND4ABX3 U14827 ( .A(n13990), .B(n12575), .C(n12574), .D(n13475), 
        .Z(n12593) );
  HS65_LL_NOR2X2 U14828 ( .A(n12867), .B(n13687), .Z(n13988) );
  HS65_LL_NOR4ABX2 U14829 ( .A(n13988), .B(n12893), .C(n12577), .D(n12576), 
        .Z(n12580) );
  HS65_LL_NOR3X1 U14830 ( .A(sa00[6]), .B(sa00[1]), .C(n12578), .Z(n13496) );
  HS65_LL_NOR4ABX2 U14831 ( .A(n12580), .B(n12579), .C(n13677), .D(n13496), 
        .Z(n14098) );
  HS65_LL_NAND4ABX3 U14832 ( .A(n14104), .B(n12582), .C(n14098), .D(n12581), 
        .Z(n12590) );
  HS65_LL_NOR2AX3 U14833 ( .A(n13684), .B(n14003), .Z(n13987) );
  HS65_LL_IVX2 U14834 ( .A(n12874), .Z(n14113) );
  HS65_LL_IVX2 U14835 ( .A(n13481), .Z(n13495) );
  HS65_LL_NAND3X2 U14836 ( .A(n13466), .B(n13487), .C(n13495), .Z(n13676) );
  HS65_LL_NOR4ABX2 U14837 ( .A(n13987), .B(n14113), .C(n12583), .D(n13676), 
        .Z(n12589) );
  HS65_LL_AOI12X2 U14838 ( .A(n12586), .B(n12585), .C(n12584), .Z(n13679) );
  HS65_LL_NAND2X2 U14839 ( .A(n13679), .B(n12587), .Z(n13501) );
  HS65_LL_NOR4ABX2 U14840 ( .A(n12589), .B(n12588), .C(n13472), .D(n13501), 
        .Z(n12898) );
  HS65_LL_NOR2X2 U14841 ( .A(n13497), .B(n14025), .Z(n14014) );
  HS65_LL_NAND4ABX3 U14842 ( .A(n12591), .B(n12590), .C(n12898), .D(n14014), 
        .Z(n12592) );
  HS65_LL_MX41X4 U14843 ( .D0(n12595), .S0(n13709), .D1(n12594), .S1(n14130), 
        .D2(n12593), .S2(n14008), .D3(n12592), .S3(n14137), .Z(n15524) );
  HS65_LL_NAND2X2 U14844 ( .A(n13517), .B(n12596), .Z(n12599) );
  HS65_LL_NOR4ABX2 U14845 ( .A(n13637), .B(n12599), .C(n12598), .D(n12597), 
        .Z(n12602) );
  HS65_LL_IVX2 U14846 ( .A(n13621), .Z(n13530) );
  HS65_LL_NOR4ABX2 U14847 ( .A(n14028), .B(n12600), .C(n13530), .D(n14053), 
        .Z(n14038) );
  HS65_LL_NOR4ABX2 U14848 ( .A(n14038), .B(n14051), .C(n13639), .D(n12616), 
        .Z(n12601) );
  HS65_LL_NAND4ABX3 U14849 ( .A(n12603), .B(n13524), .C(n12602), .D(n12601), 
        .Z(n12637) );
  HS65_LL_NAND4ABX3 U14850 ( .A(n12606), .B(n12605), .C(n12604), .D(n13506), 
        .Z(n13636) );
  HS65_LL_NAND2AX4 U14851 ( .A(n13537), .B(n12607), .Z(n13638) );
  HS65_LL_NOR4ABX2 U14852 ( .A(n12608), .B(n14041), .C(n13636), .D(n13638), 
        .Z(n12609) );
  HS65_LL_NAND4ABX3 U14853 ( .A(n13525), .B(n12616), .C(n12610), .D(n12609), 
        .Z(n12636) );
  HS65_LL_NOR2X2 U14854 ( .A(n12611), .B(n14039), .Z(n12633) );
  HS65_LL_NAND3X2 U14855 ( .A(n12613), .B(n12612), .C(n13626), .Z(n12614) );
  HS65_LL_NOR4ABX2 U14856 ( .A(n14064), .B(n12615), .C(n12633), .D(n12614), 
        .Z(n12618) );
  HS65_LL_NOR4ABX2 U14857 ( .A(n12618), .B(n12617), .C(n13553), .D(n12616), 
        .Z(n12619) );
  HS65_LL_NAND4ABX3 U14858 ( .A(n13650), .B(n13628), .C(n12620), .D(n12619), 
        .Z(n12635) );
  HS65_LL_IVX2 U14859 ( .A(n13520), .Z(n12623) );
  HS65_LL_NAND2AX4 U14860 ( .A(n12621), .B(n13511), .Z(n13536) );
  HS65_LL_NAND4ABX3 U14861 ( .A(n12623), .B(n13536), .C(n12622), .D(n14051), 
        .Z(n13635) );
  HS65_LL_AOI112X2 U14862 ( .A(sa33[5]), .B(n12625), .C(n12624), .D(n13635), 
        .Z(n12627) );
  HS65_LL_NAND3X2 U14863 ( .A(n12627), .B(n13527), .C(n12626), .Z(n12628) );
  HS65_LL_NOR3X1 U14864 ( .A(n13650), .B(n12629), .C(n12628), .Z(n14081) );
  HS65_LL_NOR4ABX2 U14865 ( .A(n14081), .B(n13621), .C(n14054), .D(n12630), 
        .Z(n12631) );
  HS65_LL_NAND4ABX3 U14866 ( .A(n12633), .B(n12632), .C(n13521), .D(n12631), 
        .Z(n12634) );
  HS65_LL_MX41X4 U14867 ( .D0(n12637), .S0(n13659), .D1(n12636), .S1(n13657), 
        .D2(n12635), .S2(n14067), .D3(n12634), .S3(n14075), .Z(n15540) );
  HS65_LLS_XOR2X3 U14868 ( .A(n15524), .B(n15540), .Z(n14089) );
  HS65_LL_OAI21X2 U14869 ( .A(n14089), .B(n12641), .C(n14808), .Z(n12640) );
  HS65_LL_IVX2 U14870 ( .A(text_in_r[116]), .Z(n12638) );
  HS65_LL_OAI212X3 U14871 ( .A(w0[20]), .B(text_in_r[116]), .C(n15255), .D(
        n12638), .E(ld_r), .Z(n12639) );
  HS65_LL_CBI4I1X3 U14872 ( .A(n12641), .B(n14089), .C(n12640), .D(n12639), 
        .Z(N262) );
  HS65_LL_NAND2X2 U14873 ( .A(n13220), .B(n14257), .Z(n13816) );
  HS65_LL_IVX2 U14874 ( .A(n12642), .Z(n12676) );
  HS65_LL_AO112X4 U14875 ( .A(n12644), .B(n12676), .C(n12643), .D(n13840), .Z(
        n12645) );
  HS65_LL_NOR4ABX2 U14876 ( .A(n12646), .B(n13210), .C(n13816), .D(n12645), 
        .Z(n14268) );
  HS65_LL_IVX2 U14877 ( .A(n12647), .Z(n13203) );
  HS65_LL_IVX2 U14878 ( .A(n13879), .Z(n13810) );
  HS65_LL_NAND3X2 U14879 ( .A(n14243), .B(n12648), .C(n13810), .Z(n12669) );
  HS65_LL_NOR3X1 U14880 ( .A(n13203), .B(n12649), .C(n12669), .Z(n13226) );
  HS65_LL_IVX2 U14881 ( .A(n12650), .Z(n13808) );
  HS65_LL_NOR3X1 U14882 ( .A(n13808), .B(n14162), .C(n14183), .Z(n12657) );
  HS65_LL_NOR2X2 U14883 ( .A(n13867), .B(n13234), .Z(n12686) );
  HS65_LL_NOR2AX3 U14884 ( .A(n14240), .B(n14161), .Z(n13814) );
  HS65_LL_NOR2X2 U14885 ( .A(n13839), .B(n14270), .Z(n13863) );
  HS65_LL_NAND3X2 U14886 ( .A(n13863), .B(n12652), .C(n12651), .Z(n12653) );
  HS65_LL_NOR4ABX2 U14887 ( .A(n12666), .B(n13814), .C(n12654), .D(n12653), 
        .Z(n14149) );
  HS65_LL_NAND3X2 U14888 ( .A(n12686), .B(n12655), .C(n14149), .Z(n12672) );
  HS65_LL_NOR4ABX2 U14889 ( .A(n12657), .B(n12656), .C(n13820), .D(n12672), 
        .Z(n12658) );
  HS65_LL_NAND3X2 U14890 ( .A(n14268), .B(n13226), .C(n12658), .Z(n12693) );
  HS65_LL_NAND3X2 U14891 ( .A(sa21[6]), .B(sa21[1]), .C(n12659), .Z(n13201) );
  HS65_LL_IVX2 U14892 ( .A(n13237), .Z(n13216) );
  HS65_LL_NOR4ABX2 U14893 ( .A(n12661), .B(n13201), .C(n13216), .D(n12660), 
        .Z(n12662) );
  HS65_LL_NAND4ABX3 U14894 ( .A(n14242), .B(n12663), .C(n12662), .D(n14157), 
        .Z(n13886) );
  HS65_LL_NAND2X2 U14895 ( .A(n12664), .B(n13841), .Z(n13832) );
  HS65_LL_NOR3X1 U14896 ( .A(n12665), .B(n14246), .C(n13832), .Z(n14147) );
  HS65_LL_IVX2 U14897 ( .A(n13210), .Z(n14165) );
  HS65_LL_NOR2X2 U14898 ( .A(n14165), .B(n14177), .Z(n13842) );
  HS65_LL_IVX2 U14899 ( .A(n14253), .Z(n14163) );
  HS65_LL_NOR4ABX2 U14900 ( .A(n12666), .B(n13842), .C(n13840), .D(n14163), 
        .Z(n12667) );
  HS65_LL_NAND4ABX3 U14901 ( .A(n12668), .B(n13886), .C(n14147), .D(n12667), 
        .Z(n12692) );
  HS65_LL_IVX2 U14902 ( .A(n14179), .Z(n14143) );
  HS65_LL_NOR4X4 U14903 ( .A(n12689), .B(n13224), .C(n12669), .D(n13882), .Z(
        n12671) );
  HS65_LL_NAND4ABX3 U14904 ( .A(n12672), .B(n14143), .C(n12671), .D(n12670), 
        .Z(n12691) );
  HS65_LL_NOR2AX3 U14905 ( .A(n13887), .B(n12673), .Z(n14264) );
  HS65_LL_OAI21X2 U14906 ( .A(n12675), .B(n12674), .C(n14264), .Z(n12688) );
  HS65_LL_AOI12X2 U14907 ( .A(n12677), .B(n12676), .C(n14183), .Z(n12685) );
  HS65_LL_NOR2X2 U14908 ( .A(n13835), .B(n13839), .Z(n13884) );
  HS65_LL_IVX2 U14909 ( .A(n12678), .Z(n14274) );
  HS65_LL_NOR3AX2 U14910 ( .A(n12680), .B(n12679), .C(n14274), .Z(n12681) );
  HS65_LL_NAND3X2 U14911 ( .A(n12682), .B(n13884), .C(n12681), .Z(n13872) );
  HS65_LL_NOR4ABX2 U14912 ( .A(n12685), .B(n12684), .C(n12683), .D(n13872), 
        .Z(n14251) );
  HS65_LL_NOR4ABX2 U14913 ( .A(n12686), .B(n13231), .C(n14165), .D(n13816), 
        .Z(n12687) );
  HS65_LL_NAND4ABX3 U14914 ( .A(n12689), .B(n12688), .C(n14251), .D(n12687), 
        .Z(n12690) );
  HS65_LL_MX41X4 U14915 ( .D0(n12693), .S0(n14283), .D1(n12692), .S1(n14285), 
        .D2(n12691), .S2(n14281), .D3(n12690), .S3(n14279), .Z(n15672) );
  HS65_LL_IVX2 U14916 ( .A(n15672), .Z(n15720) );
  HS65_LL_MUXI21X2 U14917 ( .D0(n15672), .D1(n15720), .S0(n15518), .Z(n14637)
         );
  HS65_LL_NOR2AX3 U14918 ( .A(n14575), .B(n12694), .Z(n14931) );
  HS65_LL_NAND2X2 U14919 ( .A(n14931), .B(n14587), .Z(n13125) );
  HS65_LL_NAND2X2 U14920 ( .A(n13106), .B(n13104), .Z(n15228) );
  HS65_LL_OAI21X2 U14921 ( .A(n14925), .B(n13119), .C(n15228), .Z(n14902) );
  HS65_LL_AOI12X2 U14922 ( .A(n12714), .B(n12695), .C(n14902), .Z(n12701) );
  HS65_LL_NAND2X2 U14923 ( .A(n12697), .B(n12696), .Z(n12698) );
  HS65_LL_NOR4ABX2 U14924 ( .A(n13792), .B(n12698), .C(n14573), .D(n12719), 
        .Z(n12700) );
  HS65_LL_NOR4ABX2 U14925 ( .A(n12701), .B(n12700), .C(n12699), .D(n15199), 
        .Z(n14911) );
  HS65_LL_NAND2X2 U14926 ( .A(n14911), .B(n14577), .Z(n13789) );
  HS65_LL_IVX2 U14927 ( .A(n14593), .Z(n12707) );
  HS65_LL_NAND2X2 U14928 ( .A(n14585), .B(n14584), .Z(n12704) );
  HS65_LL_NOR4ABX2 U14929 ( .A(n12705), .B(n12704), .C(n12703), .D(n12702), 
        .Z(n12706) );
  HS65_LL_NAND4ABX3 U14930 ( .A(n13798), .B(n13789), .C(n12707), .D(n12706), 
        .Z(n12748) );
  HS65_LL_NAND3X2 U14931 ( .A(n13781), .B(n12708), .C(n13785), .Z(n12709) );
  HS65_LL_NOR3X1 U14932 ( .A(n14908), .B(n12710), .C(n12709), .Z(n14598) );
  HS65_LL_AOI12X2 U14933 ( .A(n12712), .B(n13106), .C(n12711), .Z(n14915) );
  HS65_LL_NAND2X2 U14934 ( .A(n12714), .B(n12713), .Z(n13791) );
  HS65_LL_NAND3AX3 U14935 ( .A(n14903), .B(n14577), .C(n13791), .Z(n15223) );
  HS65_LL_NOR4ABX2 U14936 ( .A(n14915), .B(n13792), .C(n12715), .D(n15223), 
        .Z(n12724) );
  HS65_LL_NOR2X2 U14937 ( .A(n14922), .B(n14902), .Z(n14568) );
  HS65_LL_NAND2X2 U14938 ( .A(n12741), .B(n12716), .Z(n14590) );
  HS65_LL_NOR4ABX2 U14939 ( .A(n14568), .B(n12717), .C(n14917), .D(n14590), 
        .Z(n12718) );
  HS65_LL_NAND3X2 U14940 ( .A(n12718), .B(n14905), .C(n14601), .Z(n13126) );
  HS65_LL_NOR4ABX2 U14941 ( .A(n12721), .B(n12720), .C(n13113), .D(n12719), 
        .Z(n12723) );
  HS65_LL_NAND3X2 U14942 ( .A(n12723), .B(n12722), .C(n13096), .Z(n14927) );
  HS65_LL_NOR4ABX2 U14943 ( .A(n14598), .B(n12724), .C(n13126), .D(n14927), 
        .Z(n12746) );
  HS65_LL_IVX2 U14944 ( .A(n15238), .Z(n14935) );
  HS65_LL_OAI112X1 U14945 ( .A(n14925), .B(n12726), .C(n12725), .D(n13772), 
        .Z(n12729) );
  HS65_LL_NAND4ABX3 U14946 ( .A(n14566), .B(n12729), .C(n12728), .D(n12727), 
        .Z(n13793) );
  HS65_LL_NAND3AX3 U14947 ( .A(n12731), .B(n13100), .C(n12730), .Z(n15197) );
  HS65_LL_NAND2X2 U14948 ( .A(n14607), .B(n14580), .Z(n13121) );
  HS65_LL_NAND2AX4 U14949 ( .A(n13099), .B(n12732), .Z(n13765) );
  HS65_LL_NOR3X1 U14950 ( .A(n13780), .B(n13121), .C(n13765), .Z(n14909) );
  HS65_LL_NAND4ABX3 U14951 ( .A(n14903), .B(n15197), .C(n14909), .D(n14571), 
        .Z(n12733) );
  HS65_LL_OAI13X1 U14952 ( .A(n13793), .B(n13126), .C(n12733), .D(n15234), .Z(
        n12745) );
  HS65_LL_NOR2AX3 U14953 ( .A(n13096), .B(n13095), .Z(n12735) );
  HS65_LL_NAND4ABX3 U14954 ( .A(n13784), .B(n12736), .C(n12735), .D(n12734), 
        .Z(n13132) );
  HS65_LL_NAND4ABX3 U14955 ( .A(n12739), .B(n14611), .C(n12738), .D(n12737), 
        .Z(n15232) );
  HS65_LL_NOR4ABX2 U14956 ( .A(n14601), .B(n14580), .C(n12740), .D(n15209), 
        .Z(n12742) );
  HS65_LL_NAND4ABX3 U14957 ( .A(n13124), .B(n15232), .C(n12742), .D(n12741), 
        .Z(n12743) );
  HS65_LL_OAI13X1 U14958 ( .A(n15211), .B(n13132), .C(n12743), .D(n15236), .Z(
        n12744) );
  HS65_LL_OAI112X1 U14959 ( .A(n12746), .B(n14935), .C(n12745), .D(n12744), 
        .Z(n12747) );
  HS65_LL_CBI4I6X2 U14960 ( .A(n13125), .B(n12748), .C(n15240), .D(n12747), 
        .Z(n15249) );
  HS65_LL_MUXI21X2 U14961 ( .D0(n15248), .D1(w3[26]), .S0(n15249), .Z(n12749)
         );
  HS65_LLS_XOR3X2 U14962 ( .A(n14637), .B(n12749), .C(n15342), .Z(n12810) );
  HS65_LL_NAND2X2 U14963 ( .A(n14873), .B(n14198), .Z(n13926) );
  HS65_LL_NOR2X2 U14964 ( .A(n12750), .B(n13926), .Z(n14204) );
  HS65_LL_NOR2X2 U14965 ( .A(n14211), .B(n14210), .Z(n13897) );
  HS65_LL_NOR3X1 U14966 ( .A(n12752), .B(n13904), .C(n12751), .Z(n12753) );
  HS65_LL_NAND3X2 U14967 ( .A(n14204), .B(n13897), .C(n12753), .Z(n13140) );
  HS65_LL_NOR3X1 U14968 ( .A(n14889), .B(n12787), .C(n12754), .Z(n12755) );
  HS65_LL_NAND3X2 U14969 ( .A(n13152), .B(n12755), .C(n13162), .Z(n14877) );
  HS65_LL_NAND4ABX3 U14970 ( .A(n14864), .B(n13164), .C(n13912), .D(n12756), 
        .Z(n12757) );
  HS65_LL_NOR3X1 U14971 ( .A(n12759), .B(n12758), .C(n12757), .Z(n14217) );
  HS65_LL_NAND2X2 U14972 ( .A(n12760), .B(n12768), .Z(n14879) );
  HS65_LL_NOR4ABX2 U14973 ( .A(n12762), .B(n12761), .C(n13899), .D(n14879), 
        .Z(n12763) );
  HS65_LL_NAND4ABX3 U14974 ( .A(n13140), .B(n14877), .C(n14217), .D(n12763), 
        .Z(n12806) );
  HS65_LL_IVX2 U14975 ( .A(n13140), .Z(n12776) );
  HS65_LL_NAND4ABX3 U14976 ( .A(n13148), .B(n12765), .C(n13924), .D(n12764), 
        .Z(n12766) );
  HS65_LL_NOR4ABX2 U14977 ( .A(n12769), .B(n12768), .C(n12767), .D(n12766), 
        .Z(n13896) );
  HS65_LL_NAND2X2 U14978 ( .A(n12770), .B(n14867), .Z(n13150) );
  HS65_LL_NOR2X2 U14979 ( .A(n14863), .B(n13150), .Z(n13159) );
  HS65_LL_NAND2X2 U14980 ( .A(n13159), .B(n12771), .Z(n14885) );
  HS65_LL_NOR4ABX2 U14981 ( .A(n12773), .B(n12772), .C(n13903), .D(n14885), 
        .Z(n12775) );
  HS65_LL_AOI13X2 U14982 ( .A(n12776), .B(n13896), .C(n12775), .D(n12774), .Z(
        n12805) );
  HS65_LL_NOR2X2 U14983 ( .A(n12777), .B(n13899), .Z(n12792) );
  HS65_LL_NOR4ABX2 U14984 ( .A(n12792), .B(n13915), .C(n12778), .D(n14225), 
        .Z(n13142) );
  HS65_LL_NOR2X2 U14985 ( .A(n12780), .B(n12779), .Z(n14207) );
  HS65_LL_IVX2 U14986 ( .A(n12781), .Z(n12782) );
  HS65_LL_AOI12X2 U14987 ( .A(n12783), .B(n12782), .C(n13904), .Z(n14191) );
  HS65_LL_NAND4ABX3 U14988 ( .A(n14211), .B(n12784), .C(n14191), .D(n14867), 
        .Z(n12785) );
  HS65_LL_NOR4ABX2 U14989 ( .A(n13142), .B(n14207), .C(n12786), .D(n12785), 
        .Z(n12802) );
  HS65_LL_AOI13X2 U14990 ( .A(sa10[0]), .B(sa10[5]), .C(n12788), .D(n12787), 
        .Z(n13901) );
  HS65_LL_NOR4ABX2 U14991 ( .A(n13901), .B(n12789), .C(n14221), .D(n13926), 
        .Z(n12793) );
  HS65_LL_NOR4ABX2 U14992 ( .A(n12793), .B(n12792), .C(n12791), .D(n12790), 
        .Z(n14881) );
  HS65_LL_NAND2X2 U14993 ( .A(n14881), .B(n12794), .Z(n13920) );
  HS65_LL_NOR3X1 U14994 ( .A(n14211), .B(n12795), .C(n14219), .Z(n13931) );
  HS65_LL_NAND3X2 U14995 ( .A(n13931), .B(n12796), .C(n14212), .Z(n14876) );
  HS65_LL_NOR2X2 U14996 ( .A(n14872), .B(n12797), .Z(n14229) );
  HS65_LL_NAND4ABX3 U14997 ( .A(n12799), .B(n12798), .C(n14226), .D(n14229), 
        .Z(n12800) );
  HS65_LL_OAI13X1 U14998 ( .A(n13920), .B(n14876), .C(n12800), .D(n14891), .Z(
        n12801) );
  HS65_LL_CBI4I1X3 U14999 ( .A(n12803), .B(n12802), .C(n14895), .D(n12801), 
        .Z(n12804) );
  HS65_LL_AOI112X2 U15000 ( .A(n14893), .B(n12806), .C(n12805), .D(n12804), 
        .Z(n15343) );
  HS65_LL_OAI21X2 U15001 ( .A(n15343), .B(n12810), .C(n14832), .Z(n12809) );
  HS65_LL_IVX2 U15002 ( .A(text_in_r[26]), .Z(n12807) );
  HS65_LL_OAI212X3 U15003 ( .A(w3[26]), .B(text_in_r[26]), .C(n15248), .D(
        n12807), .E(n15545), .Z(n12808) );
  HS65_LL_CBI4I1X3 U15004 ( .A(n12810), .B(n15343), .C(n12809), .D(n12808), 
        .Z(N84) );
  HS65_LL_NAND4ABX3 U15005 ( .A(n12813), .B(n14664), .C(n12812), .D(n12811), 
        .Z(n12814) );
  HS65_LL_NOR4ABX2 U15006 ( .A(n12816), .B(n12829), .C(n12815), .D(n12814), 
        .Z(n12817) );
  HS65_LL_NAND4ABX3 U15007 ( .A(n12820), .B(n12819), .C(n12818), .D(n12817), 
        .Z(n12860) );
  HS65_LL_NAND4ABX3 U15008 ( .A(n12824), .B(n12823), .C(n12822), .D(n12821), 
        .Z(n12825) );
  HS65_LL_NOR4ABX2 U15009 ( .A(n12828), .B(n12827), .C(n12826), .D(n12825), 
        .Z(n12857) );
  HS65_LL_NAND4ABX3 U15010 ( .A(n12832), .B(n12831), .C(n12830), .D(n12829), 
        .Z(n12839) );
  HS65_LL_NOR4ABX2 U15011 ( .A(n12836), .B(n12835), .C(n12834), .D(n12833), 
        .Z(n12837) );
  HS65_LL_NAND4ABX3 U15012 ( .A(n12840), .B(n12839), .C(n12838), .D(n12837), 
        .Z(n12854) );
  HS65_LL_AOI13X2 U15013 ( .A(n12843), .B(n12842), .C(n12844), .D(n12841), .Z(
        n12848) );
  HS65_LL_NAND2AX4 U15014 ( .A(n12844), .B(n14659), .Z(n12847) );
  HS65_LL_NOR4ABX2 U15015 ( .A(n12848), .B(n12847), .C(n12846), .D(n12845), 
        .Z(n12852) );
  HS65_LL_AOI13X2 U15016 ( .A(n12852), .B(n12851), .C(n12850), .D(n12849), .Z(
        n12853) );
  HS65_LL_CBI4I6X2 U15017 ( .A(n12855), .B(n12854), .C(n14685), .D(n12853), 
        .Z(n12856) );
  HS65_LL_CBI4I1X3 U15018 ( .A(n12858), .B(n12857), .C(n14687), .D(n12856), 
        .Z(n12859) );
  HS65_LL_AOI12X2 U15019 ( .A(n14683), .B(n12860), .C(n12859), .Z(n15454) );
  HS65_LL_IVX2 U15020 ( .A(n15454), .Z(n15453) );
  HS65_LL_MUXI21X2 U15021 ( .D0(n15453), .D1(n15454), .S0(n14972), .Z(n12861)
         );
  HS65_LL_MUXI21X2 U15022 ( .D0(n14842), .D1(n14843), .S0(n12861), .Z(n12862)
         );
  HS65_LL_OAI21X2 U15023 ( .A(n11557), .B(text_in_r[88]), .C(n12862), .Z(
        n12863) );
  HS65_LLS_XNOR2X3 U15024 ( .A(w1[24]), .B(n12863), .Z(N210) );
  HS65_LL_OAI112X1 U15025 ( .A(sa00[1]), .B(sa00[6]), .C(n12865), .D(n12864), 
        .Z(n13688) );
  HS65_LL_AOI112X2 U15026 ( .A(sa00[7]), .B(n13668), .C(n12867), .D(n12866), 
        .Z(n12868) );
  HS65_LL_NAND4ABX3 U15027 ( .A(n13677), .B(n14094), .C(n13688), .D(n12868), 
        .Z(n13486) );
  HS65_LL_IVX2 U15028 ( .A(n12869), .Z(n12873) );
  HS65_LL_NOR3X1 U15029 ( .A(n14105), .B(n13695), .C(n12870), .Z(n13984) );
  HS65_LL_OAI112X1 U15030 ( .A(n12873), .B(n12872), .C(n13984), .D(n12871), 
        .Z(n12878) );
  HS65_LL_NOR4ABX2 U15031 ( .A(n13663), .B(n12875), .C(n13998), .D(n12874), 
        .Z(n12876) );
  HS65_LL_NAND4ABX3 U15032 ( .A(n13486), .B(n12878), .C(n12877), .D(n12876), 
        .Z(n12906) );
  HS65_LL_NOR4ABX2 U15033 ( .A(n14103), .B(n12885), .C(n12879), .D(n13700), 
        .Z(n12904) );
  HS65_LL_NOR4ABX2 U15034 ( .A(n12880), .B(n13488), .C(n14025), .D(n14100), 
        .Z(n12881) );
  HS65_LL_NAND3X2 U15035 ( .A(n12883), .B(n12882), .C(n12881), .Z(n14121) );
  HS65_LL_NOR4ABX2 U15036 ( .A(n12884), .B(n13490), .C(n14132), .D(n14121), 
        .Z(n12903) );
  HS65_LL_IVX2 U15037 ( .A(n12885), .Z(n12887) );
  HS65_LL_NOR4ABX2 U15038 ( .A(n13499), .B(n12888), .C(n12887), .D(n12886), 
        .Z(n12889) );
  HS65_LL_NAND4ABX3 U15039 ( .A(n12891), .B(n13695), .C(n12890), .D(n12889), 
        .Z(n12901) );
  HS65_LL_NOR4ABX2 U15040 ( .A(n12893), .B(n13986), .C(n13687), .D(n12892), 
        .Z(n12899) );
  HS65_LL_NAND3X2 U15041 ( .A(n12895), .B(n12894), .C(n13995), .Z(n13674) );
  HS65_LL_NOR4ABX2 U15042 ( .A(n12896), .B(n13488), .C(n14097), .D(n13674), 
        .Z(n12897) );
  HS65_LL_AOI13X2 U15043 ( .A(n12899), .B(n12898), .C(n12897), .D(n14134), .Z(
        n12900) );
  HS65_LL_CBI4I6X2 U15044 ( .A(n13471), .B(n12901), .C(n14137), .D(n12900), 
        .Z(n12902) );
  HS65_LL_CBI4I1X3 U15045 ( .A(n12904), .B(n12903), .C(n14125), .D(n12902), 
        .Z(n12905) );
  HS65_LL_CBI4I6X2 U15046 ( .A(n13492), .B(n12906), .C(n14130), .D(n12905), 
        .Z(n15115) );
  HS65_LL_NOR4ABX2 U15047 ( .A(n12909), .B(n12914), .C(n12908), .D(n12907), 
        .Z(n12910) );
  HS65_LL_NAND4ABX3 U15048 ( .A(n12913), .B(n12912), .C(n12911), .D(n12910), 
        .Z(n12952) );
  HS65_LL_NAND4ABX3 U15049 ( .A(n12917), .B(n12916), .C(n12915), .D(n12914), 
        .Z(n12918) );
  HS65_LL_NOR4ABX2 U15050 ( .A(n12920), .B(n12919), .C(n12928), .D(n12918), 
        .Z(n12948) );
  HS65_LL_CBI4I6X2 U15051 ( .A(n12930), .B(n12923), .C(n12922), .D(n12921), 
        .Z(n12924) );
  HS65_LL_NAND4ABX3 U15052 ( .A(n12927), .B(n12926), .C(n12925), .D(n12924), 
        .Z(n12933) );
  HS65_LL_AOI12X2 U15053 ( .A(n12930), .B(n12929), .C(n12928), .Z(n12931) );
  HS65_LL_NAND4ABX3 U15054 ( .A(n12934), .B(n12933), .C(n12932), .D(n12931), 
        .Z(n12944) );
  HS65_LL_NOR3X1 U15055 ( .A(n12937), .B(n12936), .C(n12935), .Z(n12938) );
  HS65_LL_NAND4ABX3 U15056 ( .A(n12941), .B(n12940), .C(n12939), .D(n12938), 
        .Z(n12942) );
  HS65_LL_AOI22X1 U15057 ( .A(n12945), .B(n12944), .C(n12943), .D(n12942), .Z(
        n12946) );
  HS65_LL_CBI4I1X3 U15058 ( .A(n12949), .B(n12948), .C(n12947), .D(n12946), 
        .Z(n12950) );
  HS65_LL_CBI4I6X2 U15059 ( .A(n12953), .B(n12952), .C(n12951), .D(n12950), 
        .Z(n15349) );
  HS65_LL_NAND4ABX3 U15060 ( .A(n12957), .B(n12956), .C(n12955), .D(n12954), 
        .Z(n12967) );
  HS65_LL_NAND4ABX3 U15061 ( .A(n12960), .B(n13603), .C(n12959), .D(n12958), 
        .Z(n12961) );
  HS65_LL_AOI112X2 U15062 ( .A(n12964), .B(n12963), .C(n12962), .D(n12961), 
        .Z(n12965) );
  HS65_LL_NAND4ABX3 U15063 ( .A(n12968), .B(n12967), .C(n12966), .D(n12965), 
        .Z(n13007) );
  HS65_LL_NOR4ABX2 U15064 ( .A(n12970), .B(n13573), .C(n13941), .D(n12969), 
        .Z(n12971) );
  HS65_LL_NAND4ABX3 U15065 ( .A(n12973), .B(n12972), .C(n13581), .D(n12971), 
        .Z(n13006) );
  HS65_LL_AOI112X2 U15066 ( .A(n12977), .B(n12976), .C(n12975), .D(n12974), 
        .Z(n13609) );
  HS65_LL_NOR4ABX2 U15067 ( .A(n12980), .B(n12979), .C(n13583), .D(n12978), 
        .Z(n12982) );
  HS65_LL_NOR4ABX2 U15068 ( .A(n12982), .B(n13958), .C(n12981), .D(n13950), 
        .Z(n12983) );
  HS65_LL_NAND3X2 U15069 ( .A(n12984), .B(n13609), .C(n12983), .Z(n13005) );
  HS65_LL_NOR2X2 U15070 ( .A(n12986), .B(n12985), .Z(n12995) );
  HS65_LL_NAND2AX4 U15071 ( .A(n12988), .B(n12987), .Z(n12994) );
  HS65_LL_NOR4ABX2 U15072 ( .A(n12992), .B(n12991), .C(n12990), .D(n12989), 
        .Z(n12993) );
  HS65_LL_NAND4ABX3 U15073 ( .A(n12995), .B(n12994), .C(n12993), .D(n13968), 
        .Z(n13596) );
  HS65_LL_NOR3X1 U15074 ( .A(n13942), .B(n12997), .C(n12996), .Z(n13002) );
  HS65_LL_NOR4ABX2 U15075 ( .A(n13000), .B(n13585), .C(n12999), .D(n12998), 
        .Z(n13001) );
  HS65_LL_NAND4ABX3 U15076 ( .A(n13003), .B(n13596), .C(n13002), .D(n13001), 
        .Z(n13004) );
  HS65_LL_MX41X4 U15077 ( .D0(n13007), .S0(n13961), .D1(n13006), .S1(n13972), 
        .D2(n13005), .S2(n13614), .D3(n13004), .S3(n13981), .Z(n15549) );
  HS65_LLS_XOR2X3 U15078 ( .A(n15349), .B(n15549), .Z(n15523) );
  HS65_LLS_XOR3X2 U15079 ( .A(n15115), .B(n14089), .C(n15523), .Z(n13008) );
  HS65_LL_MUXI21X2 U15080 ( .D0(n13008), .D1(text_in_r[101]), .S0(n15545), .Z(
        n13009) );
  HS65_LLS_XNOR2X3 U15081 ( .A(w0[5]), .B(n13009), .Z(N231) );
  HS65_LL_MUXI21X2 U15082 ( .D0(n15357), .D1(n15358), .S0(n14957), .Z(n13010)
         );
  HS65_LL_MUXI21X2 U15083 ( .D0(n14842), .D1(n14843), .S0(n13010), .Z(n13011)
         );
  HS65_LL_OAI21X2 U15084 ( .A(n11557), .B(text_in_r[71]), .C(n13011), .Z(
        n13012) );
  HS65_LLS_XNOR2X3 U15085 ( .A(w1[7]), .B(n13012), .Z(N169) );
  HS65_LL_OAI21X2 U15086 ( .A(w2[15]), .B(text_in_r[47]), .C(n15688), .Z(
        n13088) );
  HS65_LLS_XNOR2X3 U15087 ( .A(n15594), .B(n15277), .Z(n13013) );
  HS65_LL_NOR2AX3 U15088 ( .A(n13013), .B(n15698), .Z(n15651) );
  HS65_LL_NOR2X2 U15089 ( .A(n14822), .B(n13013), .Z(n15652) );
  HS65_LL_NOR4ABX2 U15090 ( .A(n13017), .B(n13016), .C(n13015), .D(n13014), 
        .Z(n13053) );
  HS65_LL_AOI12X2 U15091 ( .A(n13019), .B(sa20[5]), .C(n13018), .Z(n13052) );
  HS65_LL_IVX2 U15092 ( .A(n13020), .Z(n15413) );
  HS65_LL_NOR4ABX2 U15093 ( .A(n13027), .B(n13023), .C(n13022), .D(n13021), 
        .Z(n13024) );
  HS65_LL_NAND4ABX3 U15094 ( .A(n13034), .B(n13026), .C(n13025), .D(n13024), 
        .Z(n13049) );
  HS65_LL_NAND4ABX3 U15095 ( .A(n13029), .B(n13028), .C(n13027), .D(n15378), 
        .Z(n13030) );
  HS65_LL_NOR4ABX2 U15096 ( .A(n13033), .B(n13032), .C(n13031), .D(n13030), 
        .Z(n13046) );
  HS65_LL_NOR4ABX2 U15097 ( .A(n13036), .B(n13035), .C(n15407), .D(n13034), 
        .Z(n13037) );
  HS65_LL_NAND4ABX3 U15098 ( .A(n13040), .B(n13039), .C(n13038), .D(n13037), 
        .Z(n13041) );
  HS65_LL_OAI13X1 U15099 ( .A(n13043), .B(n13042), .C(n13041), .D(n15408), .Z(
        n13044) );
  HS65_LL_CBI4I1X3 U15100 ( .A(n13047), .B(n13046), .C(n13045), .D(n13044), 
        .Z(n13048) );
  HS65_LL_CBI4I6X2 U15101 ( .A(n13050), .B(n13049), .C(n15416), .D(n13048), 
        .Z(n13051) );
  HS65_LL_CBI4I1X3 U15102 ( .A(n13053), .B(n13052), .C(n15413), .D(n13051), 
        .Z(n15589) );
  HS65_LL_IVX2 U15103 ( .A(n15589), .Z(n15574) );
  HS65_LL_NOR3X1 U15104 ( .A(n13055), .B(n13080), .C(n13054), .Z(n13062) );
  HS65_LL_NOR2AX3 U15105 ( .A(n15475), .B(n13056), .Z(n13312) );
  HS65_LL_NOR4ABX2 U15106 ( .A(n13059), .B(n13312), .C(n13058), .D(n13057), 
        .Z(n13061) );
  HS65_LL_NAND3X2 U15107 ( .A(n13062), .B(n13061), .C(n13060), .Z(n13084) );
  HS65_LL_NOR3X1 U15108 ( .A(n13064), .B(n15471), .C(n13063), .Z(n15491) );
  HS65_LL_NAND4ABX3 U15109 ( .A(n13067), .B(n13066), .C(n15491), .D(n13065), 
        .Z(n13083) );
  HS65_LL_NOR2X2 U15110 ( .A(n13069), .B(n13068), .Z(n13070) );
  HS65_LL_NAND4ABX3 U15111 ( .A(n13073), .B(n13072), .C(n13071), .D(n13070), 
        .Z(n13082) );
  HS65_LL_NOR4ABX2 U15112 ( .A(n13076), .B(n13325), .C(n13075), .D(n13074), 
        .Z(n13077) );
  HS65_LL_NAND4ABX3 U15113 ( .A(n13080), .B(n13079), .C(n13078), .D(n13077), 
        .Z(n13081) );
  HS65_LL_MX41X4 U15114 ( .D0(n13084), .S0(n15478), .D1(n13083), .S1(n15494), 
        .D2(n13082), .S2(n13352), .D3(n13081), .S3(n15503), .Z(n15587) );
  HS65_LLS_XOR3X2 U15115 ( .A(n15455), .B(w2[15]), .C(n15587), .Z(n13085) );
  HS65_LL_MUXI21X2 U15116 ( .D0(n15574), .D1(n15589), .S0(n13085), .Z(n13086)
         );
  HS65_LL_MUXI21X2 U15117 ( .D0(n15651), .D1(n15652), .S0(n13086), .Z(n13087)
         );
  HS65_LL_CBI4I1X3 U15118 ( .A(text_in_r[47]), .B(w2[15]), .C(n13088), .D(
        n13087), .Z(N121) );
  HS65_LL_OAI21X2 U15119 ( .A(w2[25]), .B(text_in_r[57]), .C(n15734), .Z(
        n13093) );
  HS65_LL_MUXI21X2 U15120 ( .D0(n15426), .D1(n15425), .S0(n15511), .Z(n15608)
         );
  HS65_LL_MUXI21X2 U15121 ( .D0(n15599), .D1(n15336), .S0(w2[25]), .Z(n13089)
         );
  HS65_LLS_XOR3X2 U15122 ( .A(n15625), .B(n15608), .C(n13089), .Z(n13090) );
  HS65_LL_MUXI21X2 U15123 ( .D0(n15334), .D1(n15335), .S0(n13090), .Z(n13091)
         );
  HS65_LL_MUXI21X2 U15124 ( .D0(n15651), .D1(n15652), .S0(n13091), .Z(n13092)
         );
  HS65_LL_CBI4I1X3 U15125 ( .A(text_in_r[57]), .B(w2[25]), .C(n13093), .D(
        n13092), .Z(N147) );
  HS65_LL_OAI21X2 U15126 ( .A(w3[15]), .B(text_in_r[15]), .C(n14822), .Z(
        n13302) );
  HS65_LL_NOR4ABX2 U15127 ( .A(n13097), .B(n13096), .C(n13095), .D(n13094), 
        .Z(n13102) );
  HS65_LL_NOR4ABX2 U15128 ( .A(n13100), .B(n14580), .C(n13099), .D(n13098), 
        .Z(n13101) );
  HS65_LL_NAND4ABX3 U15129 ( .A(n13103), .B(n13794), .C(n13102), .D(n13101), 
        .Z(n13136) );
  HS65_LL_OAI21X2 U15130 ( .A(n14925), .B(n13119), .C(n13781), .Z(n14916) );
  HS65_LL_OAI21X2 U15131 ( .A(n13106), .B(n13105), .C(n13104), .Z(n14609) );
  HS65_LL_NAND3AX3 U15132 ( .A(n13108), .B(n13107), .C(n13791), .Z(n13109) );
  HS65_LL_NOR3X1 U15133 ( .A(n15215), .B(n13110), .C(n13109), .Z(n13777) );
  HS65_LL_IVX2 U15134 ( .A(n13122), .Z(n14572) );
  HS65_LL_NOR2X2 U15135 ( .A(n13766), .B(n14572), .Z(n15207) );
  HS65_LL_OAI112X1 U15136 ( .A(n13120), .B(n13111), .C(n13777), .D(n15207), 
        .Z(n13112) );
  HS65_LL_AOI112X2 U15137 ( .A(n13115), .B(n13114), .C(n13113), .D(n13112), 
        .Z(n15203) );
  HS65_LL_NOR4ABX2 U15138 ( .A(n15203), .B(n13116), .C(n14903), .D(n13127), 
        .Z(n13117) );
  HS65_LL_NAND4ABX3 U15139 ( .A(n13118), .B(n14916), .C(n14609), .D(n13117), 
        .Z(n13135) );
  HS65_LL_OAI21X2 U15140 ( .A(n13120), .B(n13119), .C(n13792), .Z(n14579) );
  HS65_LL_NOR3X1 U15141 ( .A(n14579), .B(n14596), .C(n13121), .Z(n14904) );
  HS65_LL_NOR4ABX2 U15142 ( .A(n13122), .B(n14592), .C(n15225), .D(n13765), 
        .Z(n13123) );
  HS65_LL_NAND4ABX3 U15143 ( .A(n13125), .B(n13124), .C(n14904), .D(n13123), 
        .Z(n13134) );
  HS65_LL_NAND4ABX3 U15144 ( .A(n13127), .B(n13126), .C(n13773), .D(n14924), 
        .Z(n13131) );
  HS65_LL_NOR3X1 U15145 ( .A(n13129), .B(n14573), .C(n13128), .Z(n13130) );
  HS65_LL_NAND4ABX3 U15146 ( .A(n13132), .B(n13131), .C(n13130), .D(n14592), 
        .Z(n13133) );
  HS65_LL_MX41X4 U15147 ( .D0(n13136), .S0(n15240), .D1(n13135), .S1(n15238), 
        .D2(n13134), .S2(n15236), .D3(n13133), .S3(n15234), .Z(n15194) );
  HS65_LL_AOI13X2 U15148 ( .A(sa10[7]), .B(n13138), .C(n13137), .D(n14221), 
        .Z(n13141) );
  HS65_LL_NOR4ABX2 U15149 ( .A(n13142), .B(n13141), .C(n13140), .D(n13139), 
        .Z(n13143) );
  HS65_LL_NAND3X2 U15150 ( .A(n13144), .B(n14223), .C(n13143), .Z(n13171) );
  HS65_LL_OAI21X2 U15151 ( .A(n13147), .B(n13146), .C(n13145), .Z(n13898) );
  HS65_LL_NOR4ABX2 U15152 ( .A(n13924), .B(n14190), .C(n13148), .D(n13905), 
        .Z(n13154) );
  HS65_LL_NOR4ABX2 U15153 ( .A(n13152), .B(n13151), .C(n13150), .D(n13149), 
        .Z(n13153) );
  HS65_LL_NAND4ABX3 U15154 ( .A(n13155), .B(n13898), .C(n13154), .D(n13153), 
        .Z(n13170) );
  HS65_LL_NAND2X2 U15155 ( .A(n13912), .B(n14220), .Z(n13157) );
  HS65_LL_NOR3X1 U15156 ( .A(n13899), .B(n13156), .C(n14214), .Z(n14862) );
  HS65_LL_NAND4ABX3 U15157 ( .A(n14209), .B(n13157), .C(n13931), .D(n14862), 
        .Z(n13160) );
  HS65_LL_NOR2X2 U15158 ( .A(n13906), .B(n13905), .Z(n13158) );
  HS65_LL_NAND4ABX3 U15159 ( .A(n13161), .B(n13160), .C(n13159), .D(n13158), 
        .Z(n13169) );
  HS65_LL_NAND4ABX3 U15160 ( .A(n13164), .B(n13163), .C(n14194), .D(n13162), 
        .Z(n13166) );
  HS65_LL_NOR2X2 U15161 ( .A(n13903), .B(n13926), .Z(n14866) );
  HS65_LL_NAND4ABX3 U15162 ( .A(n13167), .B(n13166), .C(n14866), .D(n13165), 
        .Z(n13168) );
  HS65_LL_MX41X4 U15163 ( .D0(n13171), .S0(n14899), .D1(n13170), .S1(n14891), 
        .D2(n13169), .S2(n14233), .D3(n13168), .S3(n14893), .Z(n15337) );
  HS65_LLS_XNOR2X3 U15164 ( .A(n15194), .B(n15337), .Z(n13172) );
  HS65_LL_NOR2AX3 U15165 ( .A(n13172), .B(n15698), .Z(n15742) );
  HS65_LL_NOR2X2 U15166 ( .A(n14822), .B(n13172), .Z(n15743) );
  HS65_LL_NAND3X2 U15167 ( .A(n13274), .B(n14720), .C(n13173), .Z(n13176) );
  HS65_LL_NOR4ABX2 U15168 ( .A(n14348), .B(n13179), .C(n14707), .D(n14376), 
        .Z(n13174) );
  HS65_LL_NAND4ABX3 U15169 ( .A(n13177), .B(n13176), .C(n13175), .D(n13174), 
        .Z(n13199) );
  HS65_LL_NAND2X2 U15170 ( .A(n13179), .B(n13178), .Z(n13268) );
  HS65_LL_IVX2 U15171 ( .A(n14371), .Z(n13262) );
  HS65_LL_NOR2X2 U15172 ( .A(n13262), .B(n13180), .Z(n13250) );
  HS65_LL_NOR4ABX2 U15173 ( .A(n13264), .B(n13260), .C(n13181), .D(n14376), 
        .Z(n13182) );
  HS65_LL_NAND4ABX3 U15174 ( .A(n13183), .B(n13268), .C(n13250), .D(n13182), 
        .Z(n13198) );
  HS65_LL_NAND4ABX3 U15175 ( .A(n14700), .B(n14718), .C(n13184), .D(n14709), 
        .Z(n13251) );
  HS65_LL_NAND4ABX3 U15176 ( .A(n13251), .B(n13185), .C(n14713), .D(n14352), 
        .Z(n13187) );
  HS65_LL_NAND4ABX3 U15177 ( .A(n13758), .B(n13187), .C(n13743), .D(n13186), 
        .Z(n13197) );
  HS65_LL_AOI12X2 U15178 ( .A(n13189), .B(n14723), .C(n13188), .Z(n13195) );
  HS65_LL_NAND4ABX3 U15179 ( .A(n13752), .B(n13191), .C(n13190), .D(n14729), 
        .Z(n13192) );
  HS65_LL_NAND4ABX3 U15180 ( .A(n14370), .B(n13192), .C(n13255), .D(n13739), 
        .Z(n13194) );
  HS65_LL_NAND4ABX3 U15181 ( .A(n13195), .B(n13194), .C(n13193), .D(n14709), 
        .Z(n13196) );
  HS65_LL_MX41X4 U15182 ( .D0(n13199), .S0(n14748), .D1(n13198), .S1(n14746), 
        .D2(n13197), .S2(n14744), .D3(n13196), .S3(n14742), .Z(n13803) );
  HS65_LL_IVX2 U15183 ( .A(n13803), .Z(n15513) );
  HS65_LL_AOI12X2 U15184 ( .A(n13200), .B(sa21[7]), .C(n14164), .Z(n14248) );
  HS65_LL_NAND2X2 U15185 ( .A(n14248), .B(n13201), .Z(n13837) );
  HS65_LL_NOR4ABX2 U15186 ( .A(n13202), .B(n14253), .C(n13232), .D(n13837), 
        .Z(n13205) );
  HS65_LL_NOR4ABX2 U15187 ( .A(n14262), .B(n13205), .C(n13204), .D(n13203), 
        .Z(n14155) );
  HS65_LL_NAND4ABX3 U15188 ( .A(n13208), .B(n13207), .C(n14155), .D(n13206), 
        .Z(n13246) );
  HS65_LL_IVX2 U15189 ( .A(n13841), .Z(n13212) );
  HS65_LL_NAND2X2 U15190 ( .A(n13210), .B(n13209), .Z(n13827) );
  HS65_LL_NOR3X1 U15191 ( .A(n13212), .B(n13211), .C(n13827), .Z(n13821) );
  HS65_LL_NOR3AX2 U15192 ( .A(n13214), .B(n13213), .C(n14177), .Z(n14275) );
  HS65_LL_NAND3X2 U15193 ( .A(n13226), .B(n13821), .C(n14275), .Z(n13219) );
  HS65_LL_NOR3X1 U15194 ( .A(n13216), .B(n14270), .C(n13215), .Z(n13217) );
  HS65_LL_NAND4ABX3 U15195 ( .A(n13872), .B(n13219), .C(n13218), .D(n13217), 
        .Z(n13245) );
  HS65_LL_NAND2X2 U15196 ( .A(n13220), .B(n14252), .Z(n14176) );
  HS65_LL_NAND4ABX3 U15197 ( .A(n13223), .B(n13222), .C(n14174), .D(n13221), 
        .Z(n13227) );
  HS65_LL_NOR2X2 U15198 ( .A(n13224), .B(n14169), .Z(n13225) );
  HS65_LL_NAND4ABX3 U15199 ( .A(n14176), .B(n13227), .C(n13226), .D(n13225), 
        .Z(n13244) );
  HS65_LL_NOR4ABX2 U15200 ( .A(n13229), .B(n13228), .C(n14144), .D(n14161), 
        .Z(n13230) );
  HS65_LL_NAND4ABX3 U15201 ( .A(n13233), .B(n13232), .C(n13231), .D(n13230), 
        .Z(n13241) );
  HS65_LL_NOR4ABX2 U15202 ( .A(n13869), .B(n13235), .C(n13234), .D(n13827), 
        .Z(n13240) );
  HS65_LL_NAND3X2 U15203 ( .A(n13237), .B(n14239), .C(n13236), .Z(n13238) );
  HS65_LL_NOR4ABX2 U15204 ( .A(n14258), .B(n13240), .C(n13239), .D(n13238), 
        .Z(n13805) );
  HS65_LL_NAND4ABX3 U15205 ( .A(n13242), .B(n13241), .C(n14271), .D(n13805), 
        .Z(n13243) );
  HS65_LL_MX41X4 U15206 ( .D0(n13246), .S0(n14285), .D1(n13245), .S1(n14283), 
        .D2(n13244), .S2(n14281), .D3(n13243), .S3(n14279), .Z(n15683) );
  HS65_LL_IVX2 U15207 ( .A(n15683), .Z(n15663) );
  HS65_LL_NOR2X2 U15208 ( .A(n13247), .B(n13740), .Z(n14365) );
  HS65_LL_NAND2X2 U15209 ( .A(n14365), .B(n13248), .Z(n13272) );
  HS65_LL_NAND4ABX3 U15210 ( .A(n13272), .B(n13251), .C(n13250), .D(n13249), 
        .Z(n13253) );
  HS65_LL_NAND4ABX3 U15211 ( .A(n13290), .B(n13253), .C(n13734), .D(n13252), 
        .Z(n13297) );
  HS65_LL_NAND3X2 U15212 ( .A(n13255), .B(n13254), .C(n14709), .Z(n14351) );
  HS65_LL_IVX2 U15213 ( .A(n14351), .Z(n14374) );
  HS65_LL_NOR3X1 U15214 ( .A(n13258), .B(n13257), .C(n13256), .Z(n13259) );
  HS65_LL_NAND3X2 U15215 ( .A(n13260), .B(n13259), .C(n14729), .Z(n13261) );
  HS65_LL_NOR4ABX2 U15216 ( .A(n14374), .B(n14720), .C(n13287), .D(n13261), 
        .Z(n14702) );
  HS65_LL_NOR4ABX2 U15217 ( .A(n13264), .B(n14702), .C(n13263), .D(n13262), 
        .Z(n13267) );
  HS65_LL_IVX2 U15218 ( .A(n14742), .Z(n13265) );
  HS65_LL_AOI13X2 U15219 ( .A(n13267), .B(n13266), .C(n14366), .D(n13265), .Z(
        n13296) );
  HS65_LL_AOI112X2 U15220 ( .A(n13271), .B(n13270), .C(n13269), .D(n13268), 
        .Z(n13273) );
  HS65_LL_NOR4ABX2 U15221 ( .A(n13274), .B(n13273), .C(n14370), .D(n13272), 
        .Z(n13755) );
  HS65_LL_NOR2X2 U15222 ( .A(n13276), .B(n13275), .Z(n13285) );
  HS65_LL_NAND2X2 U15223 ( .A(n13278), .B(n13277), .Z(n13281) );
  HS65_LL_NOR2X2 U15224 ( .A(n13287), .B(n13286), .Z(n13280) );
  HS65_LL_OAI112X1 U15225 ( .A(n13282), .B(n13281), .C(n13280), .D(n13279), 
        .Z(n13283) );
  HS65_LL_NOR4ABX2 U15226 ( .A(n13720), .B(n13285), .C(n13284), .D(n13283), 
        .Z(n13294) );
  HS65_LL_NOR3X1 U15227 ( .A(n14355), .B(n13287), .C(n13286), .Z(n14725) );
  HS65_LL_NAND4ABX3 U15228 ( .A(n13290), .B(n13289), .C(n13288), .D(n14725), 
        .Z(n13291) );
  HS65_LL_OAI13X1 U15229 ( .A(n13292), .B(n13725), .C(n13291), .D(n14746), .Z(
        n13293) );
  HS65_LL_CBI4I1X3 U15230 ( .A(n13755), .B(n13294), .C(n14380), .D(n13293), 
        .Z(n13295) );
  HS65_LL_AOI112X2 U15231 ( .A(n14748), .B(n13297), .C(n13296), .D(n13295), 
        .Z(n15682) );
  HS65_LL_MUXI21X2 U15232 ( .D0(n15683), .D1(n15663), .S0(n15682), .Z(n13298)
         );
  HS65_LL_MUXI21X2 U15233 ( .D0(n13803), .D1(n15513), .S0(n13298), .Z(n13299)
         );
  HS65_LL_MUXI21X2 U15234 ( .D0(n15427), .D1(w3[15]), .S0(n13299), .Z(n13300)
         );
  HS65_LL_MUXI21X2 U15235 ( .D0(n15742), .D1(n15743), .S0(n13300), .Z(n13301)
         );
  HS65_LL_CBI4I1X3 U15236 ( .A(text_in_r[15]), .B(w3[15]), .C(n13302), .D(
        n13301), .Z(N57) );
  HS65_LL_OAI21X2 U15237 ( .A(w2[28]), .B(text_in_r[60]), .C(n15688), .Z(
        n13359) );
  HS65_LL_IVX2 U15238 ( .A(n15419), .Z(n15420) );
  HS65_LL_AOI12X2 U15239 ( .A(n13303), .B(sa31[5]), .C(n13339), .Z(n13307) );
  HS65_LL_NOR4ABX2 U15240 ( .A(n13307), .B(n13306), .C(n13305), .D(n13304), 
        .Z(n13308) );
  HS65_LL_NAND4ABX3 U15241 ( .A(n13310), .B(n13309), .C(n13308), .D(n13317), 
        .Z(n15468) );
  HS65_LL_NOR4ABX2 U15242 ( .A(n13312), .B(n13318), .C(n13311), .D(n15468), 
        .Z(n13313) );
  HS65_LL_NAND4ABX3 U15243 ( .A(n13316), .B(n13315), .C(n13314), .D(n13313), 
        .Z(n13355) );
  HS65_LL_NAND2X2 U15244 ( .A(n13318), .B(n13317), .Z(n13323) );
  HS65_LL_NOR4ABX2 U15245 ( .A(n13319), .B(n15490), .C(n15459), .D(n13338), 
        .Z(n13320) );
  HS65_LL_NAND4ABX3 U15246 ( .A(n13323), .B(n13322), .C(n13321), .D(n13320), 
        .Z(n13354) );
  HS65_LL_IVX2 U15247 ( .A(n13324), .Z(n13326) );
  HS65_LL_NOR4ABX2 U15248 ( .A(n13326), .B(n13325), .C(n13338), .D(n15484), 
        .Z(n13333) );
  HS65_LL_NAND4ABX3 U15249 ( .A(n13329), .B(n13328), .C(n13327), .D(n15469), 
        .Z(n15480) );
  HS65_LL_NOR3X1 U15250 ( .A(n13331), .B(n15480), .C(n13330), .Z(n13332) );
  HS65_LL_NAND3X2 U15251 ( .A(n13334), .B(n13333), .C(n13332), .Z(n13353) );
  HS65_LL_NOR2X2 U15252 ( .A(n13335), .B(n15472), .Z(n13343) );
  HS65_LL_NAND4ABX3 U15253 ( .A(n13339), .B(n13338), .C(n13337), .D(n13336), 
        .Z(n13340) );
  HS65_LL_NOR4ABX2 U15254 ( .A(n13343), .B(n13342), .C(n13341), .D(n13340), 
        .Z(n13345) );
  HS65_LL_NAND4ABX3 U15255 ( .A(n13346), .B(n15462), .C(n13345), .D(n13344), 
        .Z(n13349) );
  HS65_LL_NAND4ABX3 U15256 ( .A(n13350), .B(n13349), .C(n13348), .D(n13347), 
        .Z(n13351) );
  HS65_LL_MX41X4 U15257 ( .D0(n13355), .S0(n15478), .D1(n13354), .S1(n15494), 
        .D2(n13353), .S2(n13352), .D3(n13351), .S3(n15503), .Z(n15506) );
  HS65_LL_MUXI21X2 U15258 ( .D0(n15419), .D1(n15420), .S0(n15506), .Z(n15615)
         );
  HS65_LLS_XOR3X2 U15259 ( .A(w2[28]), .B(n15615), .C(n15189), .Z(n13356) );
  HS65_LLS_XOR3X2 U15260 ( .A(n13356), .B(n15569), .C(n15331), .Z(n13357) );
  HS65_LL_MUXI21X2 U15261 ( .D0(n15651), .D1(n15652), .S0(n13357), .Z(n13358)
         );
  HS65_LL_CBI4I1X3 U15262 ( .A(text_in_r[60]), .B(w2[28]), .C(n13359), .D(
        n13358), .Z(N150) );
  HS65_LL_OAI21X2 U15263 ( .A(w2[20]), .B(text_in_r[52]), .C(n14822), .Z(
        n13364) );
  HS65_LLS_XOR2X3 U15264 ( .A(n15506), .B(n15568), .Z(n15636) );
  HS65_LL_MUXI21X2 U15265 ( .D0(n15419), .D1(n15420), .S0(w2[20]), .Z(n13360)
         );
  HS65_LLS_XOR3X2 U15266 ( .A(n15636), .B(n15579), .C(n13360), .Z(n13362) );
  HS65_LL_AOI12X2 U15267 ( .A(n13362), .B(n14627), .C(n15698), .Z(n13361) );
  HS65_LL_OAI21X2 U15268 ( .A(n13362), .B(n14627), .C(n13361), .Z(n13363) );
  HS65_LL_CBI4I1X3 U15269 ( .A(text_in_r[52]), .B(w2[20]), .C(n13364), .D(
        n13363), .Z(N134) );
  HS65_LL_OR2X4 U15270 ( .A(n13366), .B(n13365), .Z(n13374) );
  HS65_LL_NAND4ABX3 U15271 ( .A(n13370), .B(n13369), .C(n13368), .D(n13367), 
        .Z(n13373) );
  HS65_LL_NAND4ABX3 U15272 ( .A(n13374), .B(n13373), .C(n13372), .D(n13371), 
        .Z(n13411) );
  HS65_LL_NOR3X1 U15273 ( .A(n13377), .B(n13376), .C(n13375), .Z(n13380) );
  HS65_LL_NOR4ABX2 U15274 ( .A(n13381), .B(n13380), .C(n13379), .D(n13378), 
        .Z(n13385) );
  HS65_LL_NOR4ABX2 U15275 ( .A(n13385), .B(n13384), .C(n13383), .D(n13382), 
        .Z(n13408) );
  HS65_LL_NOR3X1 U15276 ( .A(n13388), .B(n13387), .C(n13386), .Z(n13389) );
  HS65_LL_OAI112X1 U15277 ( .A(n13392), .B(n13391), .C(n13390), .D(n13389), 
        .Z(n13394) );
  HS65_LL_OAI13X1 U15278 ( .A(n13396), .B(n13395), .C(n13394), .D(n13393), .Z(
        n13406) );
  HS65_LL_NAND4ABX3 U15279 ( .A(n13400), .B(n13399), .C(n13398), .D(n13397), 
        .Z(n13402) );
  HS65_LL_OAI13X1 U15280 ( .A(n13404), .B(n13403), .C(n13402), .D(n13401), .Z(
        n13405) );
  HS65_LL_OAI112X1 U15281 ( .A(n13408), .B(n13407), .C(n13406), .D(n13405), 
        .Z(n13409) );
  HS65_LL_CBI4I6X2 U15282 ( .A(n13412), .B(n13411), .C(n13410), .D(n13409), 
        .Z(n15271) );
  HS65_LL_NAND4ABX3 U15283 ( .A(n13414), .B(n13428), .C(n14320), .D(n13413), 
        .Z(n13420) );
  HS65_LL_NOR4ABX2 U15284 ( .A(n13418), .B(n13417), .C(n13416), .D(n13415), 
        .Z(n13419) );
  HS65_LL_NAND4ABX3 U15285 ( .A(n13421), .B(n13420), .C(n14300), .D(n13419), 
        .Z(n13460) );
  HS65_LL_NOR4ABX2 U15286 ( .A(n14325), .B(n13423), .C(n13422), .D(n14291), 
        .Z(n13424) );
  HS65_LL_NAND4ABX3 U15287 ( .A(n13427), .B(n13426), .C(n13425), .D(n13424), 
        .Z(n13459) );
  HS65_LL_NOR2X2 U15288 ( .A(n13429), .B(n13428), .Z(n13430) );
  HS65_LL_NAND4ABX3 U15289 ( .A(n13433), .B(n13432), .C(n13431), .D(n13430), 
        .Z(n13443) );
  HS65_LL_OAI21X2 U15290 ( .A(n13435), .B(n13434), .C(n14296), .Z(n13440) );
  HS65_LL_NAND4ABX3 U15291 ( .A(n13438), .B(n13437), .C(n13436), .D(n14325), 
        .Z(n13439) );
  HS65_LL_NOR3X1 U15292 ( .A(n13441), .B(n13440), .C(n13439), .Z(n14310) );
  HS65_LL_NAND4ABX3 U15293 ( .A(n13444), .B(n13443), .C(n14310), .D(n13442), 
        .Z(n13458) );
  HS65_LL_NOR4ABX2 U15294 ( .A(n13448), .B(n13447), .C(n13446), .D(n13445), 
        .Z(n13449) );
  HS65_LL_NAND4ABX3 U15295 ( .A(n13452), .B(n13451), .C(n13450), .D(n13449), 
        .Z(n13455) );
  HS65_LL_NAND4ABX3 U15296 ( .A(n13456), .B(n13455), .C(n13454), .D(n13453), 
        .Z(n13457) );
  HS65_LL_MX41X4 U15297 ( .D0(n13460), .S0(n14339), .D1(n13459), .S1(n14337), 
        .D2(n13458), .S2(n14335), .D3(n13457), .S3(n14333), .Z(n15365) );
  HS65_LLS_XNOR2X3 U15298 ( .A(n15271), .B(n15365), .Z(n14694) );
  HS65_LL_MUXI21X2 U15299 ( .D0(n15447), .D1(n14837), .S0(n15129), .Z(n14952)
         );
  HS65_LL_IVX2 U15300 ( .A(w1[20]), .Z(n15270) );
  HS65_LL_MUXI21X2 U15301 ( .D0(w1[20]), .D1(n15270), .S0(n15363), .Z(n13461)
         );
  HS65_LLS_XOR3X2 U15302 ( .A(n14694), .B(n14952), .C(n13461), .Z(n13465) );
  HS65_LL_OAI21X2 U15303 ( .A(n14964), .B(n13465), .C(n14832), .Z(n13464) );
  HS65_LL_IVX2 U15304 ( .A(text_in_r[84]), .Z(n13462) );
  HS65_LL_OAI212X3 U15305 ( .A(w1[20]), .B(text_in_r[84]), .C(n15270), .D(
        n13462), .E(n15545), .Z(n13463) );
  HS65_LL_CBI4I1X3 U15306 ( .A(n13465), .B(n14964), .C(n13464), .D(n13463), 
        .Z(N198) );
  HS65_LL_NAND4ABX3 U15307 ( .A(n13467), .B(n14003), .C(n14127), .D(n13466), 
        .Z(n13468) );
  HS65_LL_NOR4ABX2 U15308 ( .A(n13469), .B(n13489), .C(n14000), .D(n13468), 
        .Z(n13470) );
  HS65_LL_NAND4ABX3 U15309 ( .A(n14002), .B(n13471), .C(n14103), .D(n13470), 
        .Z(n13505) );
  HS65_LL_NAND4ABX3 U15310 ( .A(n14025), .B(n13472), .C(n14127), .D(n13487), 
        .Z(n13473) );
  HS65_LL_NAND4ABX3 U15311 ( .A(n13474), .B(n13473), .C(n13986), .D(n14114), 
        .Z(n13476) );
  HS65_LL_NAND4ABX3 U15312 ( .A(n13477), .B(n13476), .C(n14098), .D(n13475), 
        .Z(n13504) );
  HS65_LL_NOR4ABX2 U15313 ( .A(n13480), .B(n13489), .C(n13479), .D(n13478), 
        .Z(n13485) );
  HS65_LL_NOR4ABX2 U15314 ( .A(n13483), .B(n13482), .C(n13687), .D(n13481), 
        .Z(n13484) );
  HS65_LL_NAND4ABX3 U15315 ( .A(n14100), .B(n13486), .C(n13485), .D(n13484), 
        .Z(n13503) );
  HS65_LL_NAND3X2 U15316 ( .A(n13489), .B(n13488), .C(n13487), .Z(n13494) );
  HS65_LL_NAND4ABX3 U15317 ( .A(n14003), .B(n13492), .C(n13491), .D(n13490), 
        .Z(n13493) );
  HS65_LL_NOR3X1 U15318 ( .A(n13677), .B(n13494), .C(n13493), .Z(n13985) );
  HS65_LL_NAND4ABX3 U15319 ( .A(n13497), .B(n13496), .C(n13985), .D(n13495), 
        .Z(n13500) );
  HS65_LL_NAND4ABX3 U15320 ( .A(n13501), .B(n13500), .C(n13499), .D(n13498), 
        .Z(n13502) );
  HS65_LL_MX41X4 U15321 ( .D0(n13505), .S0(n13709), .D1(n13504), .S1(n14130), 
        .D2(n13503), .S2(n14008), .D3(n13502), .S3(n14137), .Z(n15553) );
  HS65_LL_NAND3X2 U15322 ( .A(n13508), .B(n13507), .C(n13506), .Z(n13509) );
  HS65_LL_NOR4ABX2 U15323 ( .A(n13512), .B(n13511), .C(n13510), .D(n13509), 
        .Z(n13513) );
  HS65_LL_NAND3X2 U15324 ( .A(n14060), .B(n13514), .C(n13513), .Z(n13563) );
  HS65_LL_AOI112X2 U15325 ( .A(n13518), .B(n13517), .C(n13516), .D(n13515), 
        .Z(n13523) );
  HS65_LL_NOR4ABX2 U15326 ( .A(n13521), .B(n13520), .C(n13519), .D(n13646), 
        .Z(n13522) );
  HS65_LL_NAND4ABX3 U15327 ( .A(n13525), .B(n13524), .C(n13523), .D(n13522), 
        .Z(n13562) );
  HS65_LL_NOR2X2 U15328 ( .A(n13630), .B(n13526), .Z(n13531) );
  HS65_LL_AND2X4 U15329 ( .A(n13528), .B(n13527), .Z(n13557) );
  HS65_LL_NOR4ABX2 U15330 ( .A(n13531), .B(n13557), .C(n13530), .D(n13529), 
        .Z(n13535) );
  HS65_LL_NOR4ABX2 U15331 ( .A(n13535), .B(n13534), .C(n13533), .D(n13532), 
        .Z(n14052) );
  HS65_LL_NOR3X1 U15332 ( .A(n13640), .B(n13537), .C(n13536), .Z(n13545) );
  HS65_LL_NAND4ABX3 U15333 ( .A(n13541), .B(n13540), .C(n13539), .D(n13538), 
        .Z(n13542) );
  HS65_LL_NOR4ABX2 U15334 ( .A(n13545), .B(n13544), .C(n13543), .D(n13542), 
        .Z(n13546) );
  HS65_LL_NAND3X2 U15335 ( .A(n13547), .B(n14052), .C(n13546), .Z(n13561) );
  HS65_LL_NAND4ABX3 U15336 ( .A(n13551), .B(n13550), .C(n13549), .D(n13548), 
        .Z(n13552) );
  HS65_LL_AOI112X2 U15337 ( .A(n13555), .B(n13554), .C(n13553), .D(n13552), 
        .Z(n13556) );
  HS65_LL_OAI112X1 U15338 ( .A(n13559), .B(n13558), .C(n13557), .D(n13556), 
        .Z(n13560) );
  HS65_LL_MX41X4 U15339 ( .D0(n13563), .S0(n13659), .D1(n13562), .S1(n13657), 
        .D2(n13561), .S2(n14067), .D3(n13560), .S3(n14075), .Z(n15551) );
  HS65_LL_IVX2 U15340 ( .A(n15551), .Z(n15550) );
  HS65_LL_MUXI21X2 U15341 ( .D0(n15550), .D1(n15551), .S0(n14633), .Z(n14793)
         );
  HS65_LLS_XOR3X2 U15342 ( .A(n15553), .B(n14793), .C(n13855), .Z(n13564) );
  HS65_LL_MUXI21X2 U15343 ( .D0(n13564), .D1(text_in_r[112]), .S0(n15545), .Z(
        n13565) );
  HS65_LLS_XNOR2X3 U15344 ( .A(w0[16]), .B(n13565), .Z(N258) );
  HS65_LL_NAND4ABX3 U15345 ( .A(n13568), .B(n13567), .C(n13607), .D(n13566), 
        .Z(n13569) );
  HS65_LL_NOR3X1 U15346 ( .A(n13571), .B(n13570), .C(n13569), .Z(n13572) );
  HS65_LL_NAND4ABX3 U15347 ( .A(n13575), .B(n13574), .C(n13573), .D(n13572), 
        .Z(n13617) );
  HS65_LL_IVX2 U15348 ( .A(n13576), .Z(n13957) );
  HS65_LL_OAI112X1 U15349 ( .A(n13579), .B(n13578), .C(n13577), .D(n13957), 
        .Z(n13580) );
  HS65_LL_NOR4ABX2 U15350 ( .A(n13582), .B(n13581), .C(n13589), .D(n13580), 
        .Z(n13584) );
  HS65_LL_NOR4ABX2 U15351 ( .A(n13607), .B(n13584), .C(n13599), .D(n13583), 
        .Z(n13586) );
  HS65_LL_NAND4ABX3 U15352 ( .A(n13588), .B(n13587), .C(n13586), .D(n13585), 
        .Z(n13616) );
  HS65_LL_AOI12X2 U15353 ( .A(n13591), .B(n13590), .C(n13589), .Z(n13595) );
  HS65_LL_NOR4ABX2 U15354 ( .A(n13949), .B(n13593), .C(n13592), .D(n13960), 
        .Z(n13594) );
  HS65_LL_NAND4ABX3 U15355 ( .A(n13597), .B(n13596), .C(n13595), .D(n13594), 
        .Z(n13615) );
  HS65_LL_NOR2X2 U15356 ( .A(n13599), .B(n13598), .Z(n13601) );
  HS65_LL_NAND4ABX3 U15357 ( .A(n13603), .B(n13602), .C(n13601), .D(n13600), 
        .Z(n13608) );
  HS65_LL_NOR2X2 U15358 ( .A(n13605), .B(n13604), .Z(n13606) );
  HS65_LL_NAND4ABX3 U15359 ( .A(n13966), .B(n13608), .C(n13607), .D(n13606), 
        .Z(n13611) );
  HS65_LL_NAND4ABX3 U15360 ( .A(n13612), .B(n13611), .C(n13610), .D(n13609), 
        .Z(n13613) );
  HS65_LL_MX41X4 U15361 ( .D0(n13617), .S0(n13961), .D1(n13616), .S1(n13972), 
        .D2(n13615), .S2(n13614), .D3(n13613), .S3(n13981), .Z(n15522) );
  HS65_LLS_XOR2X3 U15362 ( .A(n15522), .B(n15543), .Z(n14976) );
  HS65_LL_NAND3X2 U15363 ( .A(n13620), .B(n13619), .C(n13618), .Z(n14026) );
  HS65_LL_NAND3X2 U15364 ( .A(n13622), .B(n13621), .C(n13641), .Z(n13623) );
  HS65_LL_NOR3X1 U15365 ( .A(n13625), .B(n13624), .C(n13623), .Z(n13627) );
  HS65_LL_NAND4ABX3 U15366 ( .A(n13628), .B(n14026), .C(n13627), .D(n13626), 
        .Z(n13660) );
  HS65_LL_NOR4ABX2 U15367 ( .A(n13632), .B(n13631), .C(n13630), .D(n13629), 
        .Z(n13633) );
  HS65_LL_NAND4ABX3 U15368 ( .A(n13636), .B(n13635), .C(n13634), .D(n13633), 
        .Z(n13658) );
  HS65_LL_NAND4ABX3 U15369 ( .A(n13639), .B(n13638), .C(n13637), .D(n14041), 
        .Z(n13645) );
  HS65_LL_NOR4ABX2 U15370 ( .A(n13642), .B(n13641), .C(n13640), .D(n14066), 
        .Z(n13643) );
  HS65_LL_NAND4ABX3 U15371 ( .A(n13646), .B(n13645), .C(n13644), .D(n13643), 
        .Z(n13656) );
  HS65_LL_NOR3X1 U15372 ( .A(n14034), .B(n13648), .C(n13647), .Z(n13651) );
  HS65_LL_NOR4ABX2 U15373 ( .A(n14064), .B(n13651), .C(n13650), .D(n13649), 
        .Z(n13652) );
  HS65_LL_NAND3X2 U15374 ( .A(n13654), .B(n13653), .C(n13652), .Z(n13655) );
  HS65_LL_MX41X4 U15375 ( .D0(n13660), .S0(n13659), .D1(n13658), .S1(n13657), 
        .D2(n13656), .S2(n14067), .D3(n13655), .S3(n14075), .Z(n14769) );
  HS65_LL_IVX2 U15376 ( .A(n14769), .Z(n15439) );
  HS65_LL_NAND2X2 U15377 ( .A(sa00[7]), .B(n13692), .Z(n13666) );
  HS65_LL_NOR4ABX2 U15378 ( .A(n13663), .B(n13662), .C(n13661), .D(n14122), 
        .Z(n13664) );
  HS65_LL_OAI112X1 U15379 ( .A(n13666), .B(n13665), .C(n13664), .D(n14101), 
        .Z(n13667) );
  HS65_LL_AOI12X2 U15380 ( .A(sa00[1]), .B(n13668), .C(n13667), .Z(n14118) );
  HS65_LL_NAND3AX3 U15381 ( .A(n14094), .B(n13670), .C(n13669), .Z(n13671) );
  HS65_LL_NOR3X1 U15382 ( .A(n13672), .B(n14001), .C(n13671), .Z(n13673) );
  HS65_LL_NAND4ABX3 U15383 ( .A(n14010), .B(n13674), .C(n14118), .D(n13673), 
        .Z(n13710) );
  HS65_LL_NOR4ABX2 U15384 ( .A(n14013), .B(n13995), .C(n13676), .D(n13675), 
        .Z(n13678) );
  HS65_LL_NOR4ABX2 U15385 ( .A(n13679), .B(n13678), .C(n13677), .D(n14095), 
        .Z(n13680) );
  HS65_LL_NAND3X2 U15386 ( .A(n13681), .B(n13680), .C(n14101), .Z(n13708) );
  HS65_LL_NOR4ABX2 U15387 ( .A(n13685), .B(n13684), .C(n13683), .D(n13682), 
        .Z(n13690) );
  HS65_LL_NOR4ABX2 U15388 ( .A(n13688), .B(n13694), .C(n13687), .D(n13686), 
        .Z(n13689) );
  HS65_LL_NAND4ABX3 U15389 ( .A(n14121), .B(n13691), .C(n13690), .D(n13689), 
        .Z(n13707) );
  HS65_LL_NOR2X2 U15390 ( .A(n13693), .B(n13692), .Z(n13698) );
  HS65_LL_NAND2AX4 U15391 ( .A(n13695), .B(n13694), .Z(n13696) );
  HS65_LL_AOI112X2 U15392 ( .A(n13699), .B(n13698), .C(n13697), .D(n13696), 
        .Z(n13704) );
  HS65_LL_AOI112X2 U15393 ( .A(n13702), .B(sa00[1]), .C(n13701), .D(n13700), 
        .Z(n13703) );
  HS65_LL_NAND4ABX3 U15394 ( .A(n14018), .B(n13705), .C(n13704), .D(n13703), 
        .Z(n13706) );
  HS65_LL_MX41X4 U15395 ( .D0(n13710), .S0(n13709), .D1(n13708), .S1(n14130), 
        .D2(n13707), .S2(n14008), .D3(n13706), .S3(n14137), .Z(n15117) );
  HS65_LL_MUXI21X2 U15396 ( .D0(n15439), .D1(n14769), .S0(n15117), .Z(n14622)
         );
  HS65_LL_MUXI21X2 U15397 ( .D0(n15438), .D1(w0[4]), .S0(n15524), .Z(n13711)
         );
  HS65_LLS_XOR3X2 U15398 ( .A(n14976), .B(n14622), .C(n13711), .Z(n13715) );
  HS65_LLS_XOR2X3 U15399 ( .A(n15111), .B(n15435), .Z(n15556) );
  HS65_LL_OAI21X2 U15400 ( .A(n15556), .B(n13715), .C(n11557), .Z(n13714) );
  HS65_LL_IVX2 U15401 ( .A(text_in_r[100]), .Z(n13712) );
  HS65_LL_OAI212X3 U15402 ( .A(w0[4]), .B(text_in_r[100]), .C(n15438), .D(
        n13712), .E(n15545), .Z(n13713) );
  HS65_LL_CBI4I1X3 U15403 ( .A(n13715), .B(n15556), .C(n13714), .D(n13713), 
        .Z(N230) );
  HS65_LL_NAND3X2 U15404 ( .A(n13718), .B(n13717), .C(n13716), .Z(n14375) );
  HS65_LL_NAND3X2 U15405 ( .A(n13721), .B(n13720), .C(n13719), .Z(n13723) );
  HS65_LL_NAND4ABX3 U15406 ( .A(n14375), .B(n13723), .C(n14348), .D(n13722), 
        .Z(n13724) );
  HS65_LL_NOR3X1 U15407 ( .A(n13726), .B(n13725), .C(n13724), .Z(n13764) );
  HS65_LL_OAI21X2 U15408 ( .A(n13729), .B(n13728), .C(n13727), .Z(n13732) );
  HS65_LL_NOR4ABX2 U15409 ( .A(n13732), .B(n13731), .C(n13730), .D(n14370), 
        .Z(n13733) );
  HS65_LL_NAND4ABX3 U15410 ( .A(n13736), .B(n13735), .C(n13734), .D(n13733), 
        .Z(n13749) );
  HS65_LL_NOR3AX2 U15411 ( .A(n13738), .B(n13737), .C(n14707), .Z(n14349) );
  HS65_LL_NAND4ABX3 U15412 ( .A(n13741), .B(n13740), .C(n14353), .D(n13739), 
        .Z(n13742) );
  HS65_LL_NOR4ABX2 U15413 ( .A(n14349), .B(n13743), .C(n14731), .D(n13742), 
        .Z(n13745) );
  HS65_LL_AOI13X2 U15414 ( .A(n13747), .B(n13746), .C(n13745), .D(n13744), .Z(
        n13748) );
  HS65_LL_CBI4I6X2 U15415 ( .A(n13750), .B(n13749), .C(n14748), .D(n13748), 
        .Z(n13763) );
  HS65_LL_NOR3X1 U15416 ( .A(n13753), .B(n13752), .C(n13751), .Z(n13754) );
  HS65_LL_NAND3X2 U15417 ( .A(n13755), .B(n13754), .C(n14366), .Z(n14385) );
  HS65_LL_NAND4ABX3 U15418 ( .A(n13759), .B(n13758), .C(n13757), .D(n13756), 
        .Z(n13760) );
  HS65_LL_OAI13X1 U15419 ( .A(n14385), .B(n13761), .C(n13760), .D(n14742), .Z(
        n13762) );
  HS65_LL_OAI112X1 U15420 ( .A(n13764), .B(n14380), .C(n13763), .D(n13762), 
        .Z(n14760) );
  HS65_LL_IVX2 U15421 ( .A(n14760), .Z(n15516) );
  HS65_LL_NAND2X2 U15422 ( .A(n14905), .B(n14601), .Z(n13771) );
  HS65_LL_NOR4ABX2 U15423 ( .A(n13768), .B(n13767), .C(n13766), .D(n13765), 
        .Z(n13769) );
  HS65_LL_NAND4ABX3 U15424 ( .A(n14903), .B(n13771), .C(n13770), .D(n13769), 
        .Z(n13802) );
  HS65_LL_NAND3X2 U15425 ( .A(n14931), .B(n13773), .C(n13772), .Z(n13778) );
  HS65_LL_NOR4ABX2 U15426 ( .A(n14582), .B(n13775), .C(n13774), .D(n14902), 
        .Z(n13776) );
  HS65_LL_NAND4ABX3 U15427 ( .A(n15208), .B(n13778), .C(n13777), .D(n13776), 
        .Z(n13801) );
  HS65_LL_NOR2X2 U15428 ( .A(n13780), .B(n13779), .Z(n14928) );
  HS65_LL_NAND3X2 U15429 ( .A(n13782), .B(n14928), .C(n13781), .Z(n15221) );
  HS65_LL_NOR4ABX2 U15430 ( .A(n13786), .B(n13785), .C(n13784), .D(n13783), 
        .Z(n13787) );
  HS65_LL_NAND4ABX3 U15431 ( .A(n15221), .B(n13789), .C(n13788), .D(n13787), 
        .Z(n13800) );
  HS65_LL_OAI21X2 U15432 ( .A(n13790), .B(n14595), .C(n14918), .Z(n15233) );
  HS65_LL_NOR4ABX2 U15433 ( .A(n13792), .B(n13791), .C(n14590), .D(n15233), 
        .Z(n13797) );
  HS65_LL_NOR3X1 U15434 ( .A(n13795), .B(n13794), .C(n13793), .Z(n13796) );
  HS65_LL_NAND4ABX3 U15435 ( .A(n13798), .B(n14940), .C(n13797), .D(n13796), 
        .Z(n13799) );
  HS65_LL_MX41X4 U15436 ( .D0(n13802), .S0(n15240), .D1(n13801), .S1(n15238), 
        .D2(n13800), .S2(n15236), .D3(n13799), .S3(n15234), .Z(n15245) );
  HS65_LL_MUXI21X2 U15437 ( .D0(n15516), .D1(n14760), .S0(n15245), .Z(n14638)
         );
  HS65_LL_MUXI21X2 U15438 ( .D0(n15515), .D1(w3[4]), .S0(n15243), .Z(n13804)
         );
  HS65_LL_MUXI21X2 U15439 ( .D0(n13803), .D1(n15513), .S0(n15194), .Z(n15713)
         );
  HS65_LLS_XOR3X2 U15440 ( .A(n14638), .B(n13804), .C(n15713), .Z(n13853) );
  HS65_LL_NAND3X2 U15441 ( .A(n13806), .B(n13805), .C(n14173), .Z(n13807) );
  HS65_LL_NOR3X1 U15442 ( .A(n13809), .B(n13808), .C(n13807), .Z(n13862) );
  HS65_LL_IVX2 U15443 ( .A(n13837), .Z(n13813) );
  HS65_LL_NAND2X2 U15444 ( .A(n13810), .B(n13876), .Z(n13811) );
  HS65_LL_NOR4ABX2 U15445 ( .A(n13814), .B(n13813), .C(n13812), .D(n13811), 
        .Z(n13815) );
  HS65_LL_NAND4ABX3 U15446 ( .A(n14183), .B(n13816), .C(n13862), .D(n13815), 
        .Z(n13849) );
  HS65_LL_NAND3X2 U15447 ( .A(n13818), .B(n14173), .C(n13817), .Z(n13819) );
  HS65_LL_NOR4ABX2 U15448 ( .A(n13821), .B(n14257), .C(n13820), .D(n13819), 
        .Z(n13822) );
  HS65_LL_NAND3X2 U15449 ( .A(n14149), .B(n13823), .C(n13822), .Z(n13848) );
  HS65_LL_NAND2X2 U15450 ( .A(n13824), .B(n14173), .Z(n13885) );
  HS65_LL_NOR2X2 U15451 ( .A(n13826), .B(n13825), .Z(n13830) );
  HS65_LL_NOR2AX3 U15452 ( .A(n13828), .B(n13827), .Z(n14156) );
  HS65_LL_OAI13X1 U15453 ( .A(n14152), .B(n13830), .C(n13829), .D(n14156), .Z(
        n13831) );
  HS65_LL_NOR4ABX2 U15454 ( .A(n13833), .B(n13869), .C(n13832), .D(n13831), 
        .Z(n13834) );
  HS65_LL_NAND4ABX3 U15455 ( .A(n13885), .B(n13837), .C(n14264), .D(n13834), 
        .Z(n13847) );
  HS65_LL_NOR2X2 U15456 ( .A(n13835), .B(n14160), .Z(n14263) );
  HS65_LL_NAND4ABX3 U15457 ( .A(n13838), .B(n13837), .C(n13836), .D(n14263), 
        .Z(n13844) );
  HS65_LL_NOR4ABX2 U15458 ( .A(n13842), .B(n13841), .C(n13840), .D(n13839), 
        .Z(n13843) );
  HS65_LL_NAND4ABX3 U15459 ( .A(n13845), .B(n13844), .C(n14272), .D(n13843), 
        .Z(n13846) );
  HS65_LL_MX41X4 U15460 ( .D0(n13849), .S0(n14285), .D1(n13848), .S1(n14283), 
        .D2(n13847), .S2(n14281), .D3(n13846), .S3(n14279), .Z(n15428) );
  HS65_LLS_XNOR2X3 U15461 ( .A(n15338), .B(n15428), .Z(n15678) );
  HS65_LL_OAI21X2 U15462 ( .A(n15678), .B(n13853), .C(n14832), .Z(n13852) );
  HS65_LL_IVX2 U15463 ( .A(text_in_r[4]), .Z(n13850) );
  HS65_LL_OAI212X3 U15464 ( .A(w3[4]), .B(text_in_r[4]), .C(n15515), .D(n13850), .E(n15698), .Z(n13851) );
  HS65_LL_CBI4I1X3 U15465 ( .A(n13853), .B(n15678), .C(n13852), .D(n13851), 
        .Z(N38) );
  HS65_LL_MUXI21X2 U15466 ( .D0(n15257), .D1(w0[19]), .S0(n15351), .Z(n13854)
         );
  HS65_LLS_XOR3X2 U15467 ( .A(n14140), .B(n13855), .C(n13854), .Z(n13859) );
  HS65_LL_OAI21X2 U15468 ( .A(n14622), .B(n13859), .C(n14832), .Z(n13858) );
  HS65_LL_IVX2 U15469 ( .A(text_in_r[115]), .Z(n13856) );
  HS65_LL_OAI212X3 U15470 ( .A(w0[19]), .B(text_in_r[115]), .C(n15257), .D(
        n13856), .E(ld_r), .Z(n13857) );
  HS65_LL_CBI4I1X3 U15471 ( .A(n13859), .B(n14622), .C(n13858), .D(n13857), 
        .Z(N261) );
  HS65_LL_NOR4ABX2 U15472 ( .A(n13863), .B(n13862), .C(n13861), .D(n13860), 
        .Z(n13864) );
  HS65_LL_NAND4ABX3 U15473 ( .A(n13867), .B(n13866), .C(n13865), .D(n13864), 
        .Z(n13895) );
  HS65_LL_NAND2X2 U15474 ( .A(n13869), .B(n13868), .Z(n14245) );
  HS65_LL_NOR3X1 U15475 ( .A(n13872), .B(n13871), .C(n13870), .Z(n13873) );
  HS65_LL_NAND4ABX3 U15476 ( .A(n13875), .B(n14245), .C(n13874), .D(n13873), 
        .Z(n13894) );
  HS65_LL_NAND4ABX3 U15477 ( .A(n13879), .B(n13878), .C(n13877), .D(n13876), 
        .Z(n13880) );
  HS65_LL_NOR3X1 U15478 ( .A(n13882), .B(n13881), .C(n13880), .Z(n13883) );
  HS65_LL_NAND4ABX3 U15479 ( .A(n14161), .B(n14265), .C(n13884), .D(n13883), 
        .Z(n13893) );
  HS65_LL_NOR4ABX2 U15480 ( .A(n13887), .B(n14257), .C(n13886), .D(n13885), 
        .Z(n13888) );
  HS65_LL_NAND4ABX3 U15481 ( .A(n13891), .B(n13890), .C(n13889), .D(n13888), 
        .Z(n13892) );
  HS65_LL_MX41X4 U15482 ( .D0(n13895), .S0(n14285), .D1(n13894), .S1(n14283), 
        .D2(n13893), .S2(n14281), .D3(n13892), .S3(n14279), .Z(n14826) );
  HS65_LL_NAND4ABX3 U15483 ( .A(n13899), .B(n13898), .C(n13897), .D(n13896), 
        .Z(n13902) );
  HS65_LL_NAND4ABX3 U15484 ( .A(n14901), .B(n13902), .C(n13901), .D(n13900), 
        .Z(n13935) );
  HS65_LL_NOR2X2 U15485 ( .A(n13904), .B(n13903), .Z(n13909) );
  HS65_LL_NOR4ABX2 U15486 ( .A(n13907), .B(n14861), .C(n13906), .D(n13905), 
        .Z(n13908) );
  HS65_LL_NAND4ABX3 U15487 ( .A(n13911), .B(n13910), .C(n13909), .D(n13908), 
        .Z(n13934) );
  HS65_LL_IVX2 U15488 ( .A(n13912), .Z(n14227) );
  HS65_LL_NAND2X2 U15489 ( .A(n13913), .B(n14208), .Z(n13914) );
  HS65_LL_NOR4ABX2 U15490 ( .A(n13916), .B(n13915), .C(n14227), .D(n13914), 
        .Z(n13917) );
  HS65_LL_NAND4ABX3 U15491 ( .A(n13920), .B(n13919), .C(n13918), .D(n13917), 
        .Z(n13933) );
  HS65_LL_NOR4ABX2 U15492 ( .A(n13924), .B(n13923), .C(n13922), .D(n13921), 
        .Z(n13927) );
  HS65_LL_NOR4ABX2 U15493 ( .A(n13928), .B(n13927), .C(n13926), .D(n13925), 
        .Z(n13929) );
  HS65_LL_NAND3X2 U15494 ( .A(n13931), .B(n13930), .C(n13929), .Z(n13932) );
  HS65_LL_MX41X4 U15495 ( .D0(n13935), .S0(n14899), .D1(n13934), .S1(n14891), 
        .D2(n13933), .S2(n14233), .D3(n13932), .S3(n14893), .Z(n14815) );
  HS65_LLS_XOR2X3 U15496 ( .A(n14826), .B(n14815), .Z(n14761) );
  HS65_LL_MUXI21X2 U15497 ( .D0(w3[3]), .D1(n15517), .S0(n15245), .Z(n13936)
         );
  HS65_LLS_XOR3X2 U15498 ( .A(n14761), .B(n13936), .C(n15713), .Z(n13940) );
  HS65_LL_OAI21X2 U15499 ( .A(n15674), .B(n13940), .C(n14808), .Z(n13939) );
  HS65_LL_IVX2 U15500 ( .A(text_in_r[3]), .Z(n13937) );
  HS65_LL_OAI212X3 U15501 ( .A(w3[3]), .B(text_in_r[3]), .C(n15517), .D(n13937), .E(n15734), .Z(n13938) );
  HS65_LL_CBI4I1X3 U15502 ( .A(n13940), .B(n15674), .C(n13939), .D(n13938), 
        .Z(N37) );
  HS65_LL_NOR4ABX2 U15503 ( .A(n13944), .B(n13943), .C(n13942), .D(n13941), 
        .Z(n13946) );
  HS65_LL_NAND4ABX3 U15504 ( .A(n13948), .B(n13947), .C(n13946), .D(n13945), 
        .Z(n13982) );
  HS65_LL_NOR2AX3 U15505 ( .A(n13949), .B(n13960), .Z(n13952) );
  HS65_LL_NOR4ABX2 U15506 ( .A(n13953), .B(n13952), .C(n13951), .D(n13950), 
        .Z(n13956) );
  HS65_LL_NOR4ABX2 U15507 ( .A(n13964), .B(n13956), .C(n13955), .D(n13954), 
        .Z(n13979) );
  HS65_LL_NAND4ABX3 U15508 ( .A(n13960), .B(n13959), .C(n13958), .D(n13957), 
        .Z(n13962) );
  HS65_LL_OAI21X2 U15509 ( .A(n13963), .B(n13962), .C(n13961), .Z(n13977) );
  HS65_LL_NAND4ABX3 U15510 ( .A(n13967), .B(n13966), .C(n13965), .D(n13964), 
        .Z(n13974) );
  HS65_LL_NAND4ABX3 U15511 ( .A(n13971), .B(n13970), .C(n13969), .D(n13968), 
        .Z(n13973) );
  HS65_LL_OAI13X1 U15512 ( .A(n13975), .B(n13974), .C(n13973), .D(n13972), .Z(
        n13976) );
  HS65_LL_OAI112X1 U15513 ( .A(n13979), .B(n13978), .C(n13977), .D(n13976), 
        .Z(n13980) );
  HS65_LL_CBI4I6X2 U15514 ( .A(n13983), .B(n13982), .C(n13981), .D(n13980), 
        .Z(n15254) );
  HS65_LL_NAND3X2 U15515 ( .A(n13985), .B(n13984), .C(n13997), .Z(n14024) );
  HS65_LL_NAND2X2 U15516 ( .A(n14114), .B(n13986), .Z(n13989) );
  HS65_LL_NAND4ABX3 U15517 ( .A(n13990), .B(n13989), .C(n13988), .D(n13987), 
        .Z(n13991) );
  HS65_LL_NOR4ABX2 U15518 ( .A(n13994), .B(n13993), .C(n13992), .D(n13991), 
        .Z(n14022) );
  HS65_LL_AND2X4 U15519 ( .A(n13996), .B(n13995), .Z(n14123) );
  HS65_LL_NAND4ABX3 U15520 ( .A(n13999), .B(n13998), .C(n14123), .D(n13997), 
        .Z(n14099) );
  HS65_LL_NOR2X2 U15521 ( .A(n14001), .B(n14000), .Z(n14128) );
  HS65_LL_NOR3X1 U15522 ( .A(n14004), .B(n14003), .C(n14002), .Z(n14005) );
  HS65_LL_NAND4ABX3 U15523 ( .A(n14007), .B(n14006), .C(n14128), .D(n14005), 
        .Z(n14009) );
  HS65_LL_OAI13X1 U15524 ( .A(n14099), .B(n14010), .C(n14009), .D(n14008), .Z(
        n14021) );
  HS65_LL_NOR4ABX2 U15525 ( .A(n14014), .B(n14013), .C(n14012), .D(n14011), 
        .Z(n14015) );
  HS65_LL_NAND4ABX3 U15526 ( .A(n14018), .B(n14017), .C(n14016), .D(n14015), 
        .Z(n14019) );
  HS65_LL_OAI21X2 U15527 ( .A(n14099), .B(n14019), .C(n14137), .Z(n14020) );
  HS65_LL_OAI112X1 U15528 ( .A(n14022), .B(n14134), .C(n14021), .D(n14020), 
        .Z(n14023) );
  HS65_LL_CBI4I6X2 U15529 ( .A(n14025), .B(n14024), .C(n14130), .D(n14023), 
        .Z(n15113) );
  HS65_LL_NOR4ABX2 U15530 ( .A(n14029), .B(n14028), .C(n14027), .D(n14026), 
        .Z(n14032) );
  HS65_LL_NOR4ABX2 U15531 ( .A(n14032), .B(n14031), .C(n14030), .D(n14050), 
        .Z(n14080) );
  HS65_LL_AOI112X2 U15532 ( .A(n14036), .B(n14035), .C(n14034), .D(n14033), 
        .Z(n14037) );
  HS65_LL_OAI112X1 U15533 ( .A(n14040), .B(n14039), .C(n14038), .D(n14037), 
        .Z(n14077) );
  HS65_LL_NAND4ABX3 U15534 ( .A(n14044), .B(n14043), .C(n14042), .D(n14041), 
        .Z(n14076) );
  HS65_LL_NAND4ABX3 U15535 ( .A(n14048), .B(n14047), .C(n14046), .D(n14045), 
        .Z(n14049) );
  HS65_LL_NOR4ABX2 U15536 ( .A(n14052), .B(n14051), .C(n14050), .D(n14049), 
        .Z(n14055) );
  HS65_LL_NOR4ABX2 U15537 ( .A(n14056), .B(n14055), .C(n14054), .D(n14053), 
        .Z(n14072) );
  HS65_LL_NOR2X2 U15538 ( .A(n14058), .B(n14057), .Z(n14061) );
  HS65_LL_NAND4ABX3 U15539 ( .A(n14062), .B(n14061), .C(n14060), .D(n14059), 
        .Z(n14065) );
  HS65_LL_NAND4ABX3 U15540 ( .A(n14066), .B(n14065), .C(n14064), .D(n14063), 
        .Z(n14068) );
  HS65_LL_OAI21X2 U15541 ( .A(n14069), .B(n14068), .C(n14067), .Z(n14070) );
  HS65_LL_CBI4I1X3 U15542 ( .A(n14073), .B(n14072), .C(n14071), .D(n14070), 
        .Z(n14074) );
  HS65_LL_CBI4I6X2 U15543 ( .A(n14077), .B(n14076), .C(n14075), .D(n14074), 
        .Z(n14078) );
  HS65_LL_CBI4I1X3 U15544 ( .A(n14081), .B(n14080), .C(n14079), .D(n14078), 
        .Z(n15521) );
  HS65_LLS_XNOR2X3 U15545 ( .A(n15113), .B(n15521), .Z(n14980) );
  HS65_LL_MUXI21X2 U15546 ( .D0(w0[14]), .D1(n15348), .S0(n15530), .Z(n14082)
         );
  HS65_LLS_XOR3X2 U15547 ( .A(n15254), .B(n14980), .C(n14082), .Z(n14086) );
  HS65_LL_OAI21X2 U15548 ( .A(n15349), .B(n14086), .C(n14832), .Z(n14085) );
  HS65_LL_IVX2 U15549 ( .A(text_in_r[110]), .Z(n14083) );
  HS65_LL_OAI212X3 U15550 ( .A(w0[14]), .B(text_in_r[110]), .C(n15348), .D(
        n14083), .E(n15545), .Z(n14084) );
  HS65_LL_CBI4I1X3 U15551 ( .A(n14086), .B(n15349), .C(n14085), .D(n14084), 
        .Z(N248) );
  HS65_LL_OAI21X2 U15552 ( .A(w0[12]), .B(text_in_r[108]), .C(n15727), .Z(
        n14093) );
  HS65_LL_MUXI21X2 U15553 ( .D0(n15435), .D1(n15436), .S0(n15345), .Z(n14087)
         );
  HS65_LL_NOR2AX3 U15554 ( .A(n14087), .B(n15698), .Z(n14798) );
  HS65_LL_NOR2X2 U15555 ( .A(n14822), .B(n14087), .Z(n14797) );
  HS65_LL_MUXI21X2 U15556 ( .D0(w0[12]), .D1(n15350), .S0(n15439), .Z(n14088)
         );
  HS65_LLS_XOR3X2 U15557 ( .A(n14089), .B(n15522), .C(n14088), .Z(n14090) );
  HS65_LL_MUX21I1X3 U15558 ( .D0(n15351), .D1(n15351), .S0(n14090), .Z(n14091)
         );
  HS65_LL_MUXI21X2 U15559 ( .D0(n14798), .D1(n14797), .S0(n14091), .Z(n14092)
         );
  HS65_LL_CBI4I1X3 U15560 ( .A(text_in_r[108]), .B(w0[12]), .C(n14093), .D(
        n14092), .Z(N246) );
  HS65_LL_NOR2X2 U15561 ( .A(n14095), .B(n14094), .Z(n14112) );
  HS65_LL_NOR4ABX2 U15562 ( .A(n14098), .B(n14112), .C(n14097), .D(n14096), 
        .Z(n14124) );
  HS65_LL_NOR4ABX2 U15563 ( .A(n14124), .B(n14101), .C(n14100), .D(n14099), 
        .Z(n14102) );
  HS65_LL_NAND4ABX3 U15564 ( .A(n14105), .B(n14104), .C(n14103), .D(n14102), 
        .Z(n14138) );
  HS65_LL_NAND2X2 U15565 ( .A(sa00[3]), .B(sa00[0]), .Z(n14116) );
  HS65_LL_OAI112X1 U15566 ( .A(n14108), .B(n14116), .C(n14107), .D(n14106), 
        .Z(n14109) );
  HS65_LL_NOR4ABX2 U15567 ( .A(n14112), .B(n14111), .C(n14110), .D(n14109), 
        .Z(n14135) );
  HS65_LL_OAI112X1 U15568 ( .A(n14116), .B(n14115), .C(n14114), .D(n14113), 
        .Z(n14119) );
  HS65_LL_NAND4ABX3 U15569 ( .A(n14120), .B(n14119), .C(n14118), .D(n14117), 
        .Z(n14131) );
  HS65_LL_NOR4ABX2 U15570 ( .A(n14124), .B(n14123), .C(n14122), .D(n14121), 
        .Z(n14126) );
  HS65_LL_AOI13X2 U15571 ( .A(n14128), .B(n14127), .C(n14126), .D(n14125), .Z(
        n14129) );
  HS65_LL_CBI4I6X2 U15572 ( .A(n14132), .B(n14131), .C(n14130), .D(n14129), 
        .Z(n14133) );
  HS65_LL_OAI21X2 U15573 ( .A(n14135), .B(n14134), .C(n14133), .Z(n14136) );
  HS65_LL_CBI4I6X2 U15574 ( .A(n14139), .B(n14138), .C(n14137), .D(n14136), 
        .Z(n15119) );
  HS65_LLS_XOR2X3 U15575 ( .A(n15552), .B(n15441), .Z(n14794) );
  HS65_LLS_XOR3X2 U15576 ( .A(n15119), .B(n14794), .C(n14140), .Z(n14141) );
  HS65_LL_MUXI21X2 U15577 ( .D0(n14141), .D1(text_in_r[98]), .S0(n15545), .Z(
        n14142) );
  HS65_LLS_XNOR2X3 U15578 ( .A(w0[2]), .B(n14142), .Z(N228) );
  HS65_LLS_XNOR2X3 U15579 ( .A(n15249), .B(n15519), .Z(n15719) );
  HS65_LL_MUXI21X2 U15580 ( .D0(w3[17]), .D1(n15344), .S0(n15432), .Z(n14237)
         );
  HS65_LL_NOR3X1 U15581 ( .A(n14144), .B(n14183), .C(n14143), .Z(n14146) );
  HS65_LL_NOR4ABX2 U15582 ( .A(n14147), .B(n14146), .C(n14265), .D(n14145), 
        .Z(n14148) );
  HS65_LL_NAND3X2 U15583 ( .A(n14149), .B(n14272), .C(n14148), .Z(n14187) );
  HS65_LL_AOI12X2 U15584 ( .A(n14152), .B(n14151), .C(n14150), .Z(n14159) );
  HS65_LL_NOR4ABX2 U15585 ( .A(n14156), .B(n14155), .C(n14154), .D(n14153), 
        .Z(n14158) );
  HS65_LL_NAND3X2 U15586 ( .A(n14159), .B(n14158), .C(n14157), .Z(n14186) );
  HS65_LL_NOR2X2 U15587 ( .A(n14161), .B(n14160), .Z(n14254) );
  HS65_LL_NOR2X2 U15588 ( .A(n14163), .B(n14162), .Z(n14181) );
  HS65_LL_NAND4ABX3 U15589 ( .A(n14165), .B(n14164), .C(n14254), .D(n14181), 
        .Z(n14172) );
  HS65_LL_NAND4ABX3 U15590 ( .A(n14169), .B(n14168), .C(n14167), .D(n14166), 
        .Z(n14171) );
  HS65_LL_NAND4ABX3 U15591 ( .A(n14172), .B(n14171), .C(n14272), .D(n14170), 
        .Z(n14185) );
  HS65_LL_NAND3X2 U15592 ( .A(n14175), .B(n14174), .C(n14173), .Z(n14182) );
  HS65_LL_NOR4ABX2 U15593 ( .A(n14179), .B(n14178), .C(n14177), .D(n14176), 
        .Z(n14180) );
  HS65_LL_NAND4ABX3 U15594 ( .A(n14183), .B(n14182), .C(n14181), .D(n14180), 
        .Z(n14184) );
  HS65_LL_MX41X4 U15595 ( .D0(n14187), .S0(n14285), .D1(n14186), .S1(n14283), 
        .D2(n14185), .S2(n14281), .D3(n14184), .S3(n14279), .Z(n15667) );
  HS65_LL_IVX2 U15596 ( .A(n15667), .Z(n15434) );
  HS65_LL_AND2X4 U15597 ( .A(n14212), .B(n14188), .Z(n14193) );
  HS65_LL_NOR4ABX2 U15598 ( .A(n14191), .B(n14190), .C(n14209), .D(n14189), 
        .Z(n14192) );
  HS65_LL_NAND3X2 U15599 ( .A(n14194), .B(n14193), .C(n14192), .Z(n14888) );
  HS65_LL_AOI112X2 U15600 ( .A(n14197), .B(n14196), .C(n14195), .D(n14888), 
        .Z(n14199) );
  HS65_LL_NAND4ABX3 U15601 ( .A(n14201), .B(n14200), .C(n14199), .D(n14198), 
        .Z(n14236) );
  HS65_LL_NAND4ABX3 U15602 ( .A(n14213), .B(n14202), .C(n14226), .D(n14215), 
        .Z(n14205) );
  HS65_LL_NAND4ABX3 U15603 ( .A(n14206), .B(n14205), .C(n14204), .D(n14203), 
        .Z(n14235) );
  HS65_LL_NAND4ABX3 U15604 ( .A(n14210), .B(n14209), .C(n14208), .D(n14207), 
        .Z(n14218) );
  HS65_LL_NOR2AX3 U15605 ( .A(n14212), .B(n14211), .Z(n14880) );
  HS65_LL_NOR4ABX2 U15606 ( .A(n14215), .B(n14880), .C(n14214), .D(n14213), 
        .Z(n14216) );
  HS65_LL_NAND4ABX3 U15607 ( .A(n14219), .B(n14218), .C(n14217), .D(n14216), 
        .Z(n14234) );
  HS65_LL_NAND2AX4 U15608 ( .A(n14221), .B(n14220), .Z(n14224) );
  HS65_LL_NAND4ABX3 U15609 ( .A(n14225), .B(n14224), .C(n14223), .D(n14222), 
        .Z(n14231) );
  HS65_LL_NAND4ABX3 U15610 ( .A(n14227), .B(n14879), .C(n14226), .D(n14867), 
        .Z(n14230) );
  HS65_LL_NAND4ABX3 U15611 ( .A(n14231), .B(n14230), .C(n14229), .D(n14228), 
        .Z(n14232) );
  HS65_LL_MX41X4 U15612 ( .D0(n14236), .S0(n14899), .D1(n14235), .S1(n14891), 
        .D2(n14234), .S2(n14233), .D3(n14232), .S3(n14893), .Z(n15693) );
  HS65_LL_MUXI21X2 U15613 ( .D0(n15667), .D1(n15434), .S0(n15693), .Z(n15712)
         );
  HS65_LLS_XOR3X2 U15614 ( .A(n15719), .B(n14237), .C(n15712), .Z(n14290) );
  HS65_LL_NAND3X2 U15615 ( .A(n14240), .B(n14239), .C(n14238), .Z(n14241) );
  HS65_LL_NOR4ABX2 U15616 ( .A(n14244), .B(n14243), .C(n14242), .D(n14241), 
        .Z(n14250) );
  HS65_LL_NOR4ABX2 U15617 ( .A(n14248), .B(n14247), .C(n14246), .D(n14245), 
        .Z(n14249) );
  HS65_LL_NAND3X2 U15618 ( .A(n14251), .B(n14250), .C(n14249), .Z(n14286) );
  HS65_LL_NAND3X2 U15619 ( .A(n14254), .B(n14253), .C(n14252), .Z(n14260) );
  HS65_LL_NOR4ABX2 U15620 ( .A(n14258), .B(n14257), .C(n14256), .D(n14255), 
        .Z(n14259) );
  HS65_LL_NAND4ABX3 U15621 ( .A(n14261), .B(n14260), .C(n14264), .D(n14259), 
        .Z(n14284) );
  HS65_LL_NAND3X2 U15622 ( .A(n14264), .B(n14263), .C(n14262), .Z(n14269) );
  HS65_LL_AOI13X2 U15623 ( .A(sa21[5]), .B(sa21[3]), .C(n14266), .D(n14265), 
        .Z(n14267) );
  HS65_LL_NAND4ABX3 U15624 ( .A(n14270), .B(n14269), .C(n14268), .D(n14267), 
        .Z(n14282) );
  HS65_LL_NAND4ABX3 U15625 ( .A(n14274), .B(n14273), .C(n14272), .D(n14271), 
        .Z(n14277) );
  HS65_LL_NAND4ABX3 U15626 ( .A(n14278), .B(n14277), .C(n14276), .D(n14275), 
        .Z(n14280) );
  HS65_LL_MX41X4 U15627 ( .D0(n14286), .S0(n14285), .D1(n14284), .S1(n14283), 
        .D2(n14282), .S2(n14281), .D3(n14280), .S3(n14279), .Z(n15740) );
  HS65_LL_IVX2 U15628 ( .A(n15740), .Z(n15739) );
  HS65_LL_MUXI21X2 U15629 ( .D0(n15739), .D1(n15740), .S0(n15337), .Z(n15668)
         );
  HS65_LL_OAI21X2 U15630 ( .A(n15668), .B(n14290), .C(n14832), .Z(n14289) );
  HS65_LL_IVX2 U15631 ( .A(text_in_r[17]), .Z(n14287) );
  HS65_LL_OAI212X3 U15632 ( .A(w3[17]), .B(text_in_r[17]), .C(n15344), .D(
        n14287), .E(n15545), .Z(n14288) );
  HS65_LL_CBI4I1X3 U15633 ( .A(n14290), .B(n15668), .C(n14289), .D(n14288), 
        .Z(N67) );
  HS65_LL_NOR2X2 U15634 ( .A(n14292), .B(n14291), .Z(n14321) );
  HS65_LL_NAND4ABX3 U15635 ( .A(n14295), .B(n14294), .C(n14293), .D(n14321), 
        .Z(n14327) );
  HS65_LL_NAND2X2 U15636 ( .A(n14297), .B(n14296), .Z(n14303) );
  HS65_LL_NOR4ABX2 U15637 ( .A(n14300), .B(n14314), .C(n14299), .D(n14298), 
        .Z(n14301) );
  HS65_LL_NAND4ABX3 U15638 ( .A(n14327), .B(n14303), .C(n14302), .D(n14301), 
        .Z(n14340) );
  HS65_LL_AOI12X2 U15639 ( .A(n14306), .B(n14305), .C(n14304), .Z(n14308) );
  HS65_LL_OAI112X1 U15640 ( .A(n14309), .B(n14316), .C(n14308), .D(n14307), 
        .Z(n14312) );
  HS65_LL_NAND4ABX3 U15641 ( .A(n14313), .B(n14312), .C(n14311), .D(n14310), 
        .Z(n14338) );
  HS65_LL_OAI112X1 U15642 ( .A(n14317), .B(n14316), .C(n14315), .D(n14314), 
        .Z(n14318) );
  HS65_LL_NOR4ABX2 U15643 ( .A(n14321), .B(n14320), .C(n14319), .D(n14318), 
        .Z(n14322) );
  HS65_LL_NAND3X2 U15644 ( .A(n14324), .B(n14323), .C(n14322), .Z(n14336) );
  HS65_LL_NAND4ABX3 U15645 ( .A(n14328), .B(n14327), .C(n14326), .D(n14325), 
        .Z(n14331) );
  HS65_LL_NAND4ABX3 U15646 ( .A(n14332), .B(n14331), .C(n14330), .D(n14329), 
        .Z(n14334) );
  HS65_LL_MX41X4 U15647 ( .D0(n14340), .S0(n14339), .D1(n14338), .S1(n14337), 
        .D2(n14336), .S2(n14335), .D3(n14334), .S3(n14333), .Z(n15367) );
  HS65_LL_IVX2 U15648 ( .A(n15367), .Z(n15368) );
  HS65_LL_MUXI21X2 U15649 ( .D0(n15367), .D1(n15368), .S0(n14647), .Z(n14778)
         );
  HS65_LL_IVX2 U15650 ( .A(w1[26]), .Z(n15134) );
  HS65_LL_MUXI21X2 U15651 ( .D0(w1[26]), .D1(n15134), .S0(n15273), .Z(n14341)
         );
  HS65_LLS_XOR3X2 U15652 ( .A(n14778), .B(n14341), .C(n15135), .Z(n14345) );
  HS65_LL_OAI21X2 U15653 ( .A(n14854), .B(n14345), .C(n14832), .Z(n14344) );
  HS65_LL_IVX2 U15654 ( .A(text_in_r[90]), .Z(n14342) );
  HS65_LL_OAI212X3 U15655 ( .A(w1[26]), .B(text_in_r[90]), .C(n15134), .D(
        n14342), .E(n15545), .Z(n14343) );
  HS65_LL_CBI4I1X3 U15656 ( .A(n14345), .B(n14854), .C(n14344), .D(n14343), 
        .Z(N212) );
  HS65_LL_IVX2 U15657 ( .A(n14737), .Z(n14347) );
  HS65_LL_NOR4ABX2 U15658 ( .A(n14349), .B(n14348), .C(n14347), .D(n14346), 
        .Z(n14350) );
  HS65_LL_NAND4ABX3 U15659 ( .A(n14735), .B(n14351), .C(n14350), .D(n14703), 
        .Z(n14384) );
  HS65_LL_NAND2X2 U15660 ( .A(n14352), .B(n14371), .Z(n14734) );
  HS65_LL_NAND4ABX3 U15661 ( .A(n14355), .B(n14734), .C(n14354), .D(n14353), 
        .Z(n14356) );
  HS65_LL_NOR4ABX2 U15662 ( .A(n14374), .B(n14357), .C(n14708), .D(n14356), 
        .Z(n14381) );
  HS65_LL_NOR4ABX2 U15663 ( .A(n14361), .B(n14360), .C(n14359), .D(n14358), 
        .Z(n14362) );
  HS65_LL_NAND4ABX3 U15664 ( .A(n14741), .B(n14363), .C(n14365), .D(n14362), 
        .Z(n14378) );
  HS65_LL_NAND3X2 U15665 ( .A(n14365), .B(n14364), .C(n14728), .Z(n14705) );
  HS65_LL_NAND4ABX3 U15666 ( .A(n14368), .B(n14705), .C(n14367), .D(n14366), 
        .Z(n14369) );
  HS65_LL_NOR4ABX2 U15667 ( .A(n14372), .B(n14371), .C(n14370), .D(n14369), 
        .Z(n14373) );
  HS65_LL_NAND4ABX3 U15668 ( .A(n14376), .B(n14375), .C(n14374), .D(n14373), 
        .Z(n14377) );
  HS65_LL_AOI22X1 U15669 ( .A(n14748), .B(n14378), .C(n14746), .D(n14377), .Z(
        n14379) );
  HS65_LL_CBI4I1X3 U15670 ( .A(n14382), .B(n14381), .C(n14380), .D(n14379), 
        .Z(n14383) );
  HS65_LL_CBI4I6X2 U15671 ( .A(n14385), .B(n14384), .C(n14742), .D(n14383), 
        .Z(n15514) );
  HS65_LL_IVX2 U15672 ( .A(n15514), .Z(n14823) );
  HS65_LL_MUXI21X2 U15673 ( .D0(n15514), .D1(n14823), .S0(n15428), .Z(n15704)
         );
  HS65_LL_IVX2 U15674 ( .A(w3[20]), .Z(n15339) );
  HS65_LL_MUXI21X2 U15675 ( .D0(w3[20]), .D1(n15339), .S0(n15243), .Z(n14386)
         );
  HS65_LLS_XOR3X2 U15676 ( .A(n15668), .B(n15704), .C(n14386), .Z(n14390) );
  HS65_LL_OAI21X2 U15677 ( .A(n14761), .B(n14390), .C(n14832), .Z(n14389) );
  HS65_LL_IVX2 U15678 ( .A(text_in_r[20]), .Z(n14387) );
  HS65_LL_OAI212X3 U15679 ( .A(w3[20]), .B(text_in_r[20]), .C(n15339), .D(
        n14387), .E(ld_r), .Z(n14388) );
  HS65_LL_CBI4I1X3 U15680 ( .A(n14390), .B(n14761), .C(n14389), .D(n14388), 
        .Z(N70) );
  HS65_LL_MUXI21X2 U15681 ( .D0(w3[19]), .D1(n15341), .S0(n14826), .Z(n14392)
         );
  HS65_LL_MUXI21X2 U15682 ( .D0(n15672), .D1(n15720), .S0(n15342), .Z(n14391)
         );
  HS65_LLS_XOR3X2 U15683 ( .A(n15668), .B(n14392), .C(n14391), .Z(n14396) );
  HS65_LL_OAI21X2 U15684 ( .A(n14638), .B(n14396), .C(n14808), .Z(n14395) );
  HS65_LL_IVX2 U15685 ( .A(text_in_r[19]), .Z(n14393) );
  HS65_LL_OAI212X3 U15686 ( .A(w3[19]), .B(text_in_r[19]), .C(n15341), .D(
        n14393), .E(n15698), .Z(n14394) );
  HS65_LL_CBI4I1X3 U15687 ( .A(n14396), .B(n14638), .C(n14395), .D(n14394), 
        .Z(N69) );
  HS65_LL_OAI21X2 U15688 ( .A(w2[9]), .B(text_in_r[41]), .C(n15688), .Z(n14401) );
  HS65_LLS_XNOR2X3 U15689 ( .A(n15455), .B(n15649), .Z(n14397) );
  HS65_LL_NOR2AX3 U15690 ( .A(n14397), .B(n15698), .Z(n15603) );
  HS65_LL_NOR2X2 U15691 ( .A(n14822), .B(n14397), .Z(n15602) );
  HS65_LLS_XOR3X2 U15692 ( .A(w2[9]), .B(n15561), .C(n15578), .Z(n14398) );
  HS65_LLS_XOR3X2 U15693 ( .A(n15631), .B(n14398), .C(n15334), .Z(n14399) );
  HS65_LL_MUXI21X2 U15694 ( .D0(n15603), .D1(n15602), .S0(n14399), .Z(n14400)
         );
  HS65_LL_CBI4I1X3 U15695 ( .A(text_in_r[41]), .B(w2[9]), .C(n14401), .D(
        n14400), .Z(N115) );
  HS65_LL_IVX2 U15696 ( .A(n15124), .Z(n15123) );
  HS65_LL_MUXI21X2 U15697 ( .D0(n15124), .D1(n15123), .S0(n15443), .Z(n14973)
         );
  HS65_LL_IVX2 U15698 ( .A(w1[1]), .Z(n15452) );
  HS65_LL_MUXI21X2 U15699 ( .D0(n15452), .D1(w1[1]), .S0(n15135), .Z(n14402)
         );
  HS65_LLS_XOR3X2 U15700 ( .A(n14968), .B(n14973), .C(n14402), .Z(n14406) );
  HS65_LLS_XNOR2X3 U15701 ( .A(n15454), .B(n15137), .Z(n14965) );
  HS65_LL_OAI21X2 U15702 ( .A(n14965), .B(n14406), .C(n14832), .Z(n14405) );
  HS65_LL_IVX2 U15703 ( .A(text_in_r[65]), .Z(n14403) );
  HS65_LL_OAI212X3 U15704 ( .A(w1[1]), .B(text_in_r[65]), .C(n15452), .D(
        n14403), .E(ld_r), .Z(n14404) );
  HS65_LL_CBI4I1X3 U15705 ( .A(n14406), .B(n14965), .C(n14405), .D(n14404), 
        .Z(N163) );
  HS65_LL_IVX2 U15706 ( .A(w1[3]), .Z(n15450) );
  HS65_LL_NAND4ABX3 U15707 ( .A(n14410), .B(n14409), .C(n14408), .D(n14407), 
        .Z(n14413) );
  HS65_LL_NAND4ABX3 U15708 ( .A(n14414), .B(n14413), .C(n14412), .D(n14411), 
        .Z(n14454) );
  HS65_LL_NOR4ABX2 U15709 ( .A(n14418), .B(n14417), .C(n14416), .D(n14415), 
        .Z(n14420) );
  HS65_LL_NAND4ABX3 U15710 ( .A(n14422), .B(n14421), .C(n14420), .D(n14419), 
        .Z(n14452) );
  HS65_LL_NAND2AX4 U15711 ( .A(n14424), .B(n14423), .Z(n14435) );
  HS65_LL_NOR3X1 U15712 ( .A(n14427), .B(n14426), .C(n14425), .Z(n14428) );
  HS65_LL_OAI112X1 U15713 ( .A(n14431), .B(n14430), .C(n14429), .D(n14428), 
        .Z(n14434) );
  HS65_LL_NAND4ABX3 U15714 ( .A(n14435), .B(n14434), .C(n14433), .D(n14432), 
        .Z(n14450) );
  HS65_LL_NOR3X1 U15715 ( .A(n14438), .B(n14437), .C(n14436), .Z(n14439) );
  HS65_LL_NAND4ABX3 U15716 ( .A(n14442), .B(n14441), .C(n14440), .D(n14439), 
        .Z(n14445) );
  HS65_LL_NAND4ABX3 U15717 ( .A(n14446), .B(n14445), .C(n14444), .D(n14443), 
        .Z(n14448) );
  HS65_LL_MX41X4 U15718 ( .D0(n14454), .S0(n14453), .D1(n14452), .S1(n14451), 
        .D2(n14450), .S2(n14449), .D3(n14448), .S3(n14447), .Z(n15131) );
  HS65_LL_MUXI21X2 U15719 ( .D0(n15450), .D1(w1[3]), .S0(n15131), .Z(n14455)
         );
  HS65_LLS_XOR3X2 U15720 ( .A(n14694), .B(n14973), .C(n14455), .Z(n14459) );
  HS65_LL_OAI21X2 U15721 ( .A(n14969), .B(n14459), .C(n14832), .Z(n14458) );
  HS65_LL_IVX2 U15722 ( .A(text_in_r[67]), .Z(n14456) );
  HS65_LL_OAI212X3 U15723 ( .A(w1[3]), .B(text_in_r[67]), .C(n15450), .D(
        n14456), .E(n15734), .Z(n14457) );
  HS65_LL_CBI4I1X3 U15724 ( .A(n14459), .B(n14969), .C(n14458), .D(n14457), 
        .Z(N165) );
  HS65_LL_OAI21X2 U15725 ( .A(w2[12]), .B(text_in_r[44]), .C(n15688), .Z(
        n14465) );
  HS65_LL_IVX2 U15726 ( .A(w2[12]), .Z(n14460) );
  HS65_LL_MUXI21X2 U15727 ( .D0(n14460), .D1(w2[12]), .S0(n15421), .Z(n14461)
         );
  HS65_LLS_XOR3X2 U15728 ( .A(n15636), .B(n15569), .C(n14461), .Z(n14462) );
  HS65_LL_MUXI21X2 U15729 ( .D0(n14628), .D1(n15508), .S0(n14462), .Z(n14463)
         );
  HS65_LL_MUXI21X2 U15730 ( .D0(n15602), .D1(n15603), .S0(n14463), .Z(n14464)
         );
  HS65_LL_CBI4I1X3 U15731 ( .A(text_in_r[44]), .B(w2[12]), .C(n14465), .D(
        n14464), .Z(N118) );
  HS65_LL_OAI21X2 U15732 ( .A(w2[31]), .B(text_in_r[63]), .C(n15727), .Z(
        n14541) );
  HS65_LL_NAND4ABX3 U15733 ( .A(n14469), .B(n14468), .C(n14467), .D(n14466), 
        .Z(n14472) );
  HS65_LL_NAND4ABX3 U15734 ( .A(n14483), .B(n14472), .C(n14471), .D(n14470), 
        .Z(n14500) );
  HS65_LL_IVX2 U15735 ( .A(n14473), .Z(n15151) );
  HS65_LL_NOR4ABX2 U15736 ( .A(n14476), .B(n15151), .C(n14475), .D(n14474), 
        .Z(n14479) );
  HS65_LL_NOR4ABX2 U15737 ( .A(n14480), .B(n14479), .C(n14478), .D(n14477), 
        .Z(n14481) );
  HS65_LL_NAND3AX3 U15738 ( .A(n14483), .B(n14482), .C(n14481), .Z(n14499) );
  HS65_LL_NAND3X2 U15739 ( .A(n14485), .B(n15162), .C(n14484), .Z(n14492) );
  HS65_LL_NAND4ABX3 U15740 ( .A(n14488), .B(n14487), .C(n14486), .D(n15144), 
        .Z(n14491) );
  HS65_LL_NAND4ABX3 U15741 ( .A(n14492), .B(n14491), .C(n14490), .D(n14489), 
        .Z(n14498) );
  HS65_LL_NAND4ABX3 U15742 ( .A(n14496), .B(n14495), .C(n14494), .D(n14493), 
        .Z(n14497) );
  HS65_LL_MX41X4 U15743 ( .D0(n14500), .S0(n15186), .D1(n14499), .S1(n15184), 
        .D2(n14498), .S2(n15182), .D3(n14497), .S3(n15180), .Z(n15641) );
  HS65_LL_NAND4ABX3 U15744 ( .A(n14503), .B(n14502), .C(n14530), .D(n14501), 
        .Z(n14504) );
  HS65_LL_NOR3X1 U15745 ( .A(n14506), .B(n14505), .C(n14504), .Z(n14507) );
  HS65_LL_NAND4ABX3 U15746 ( .A(n14510), .B(n14509), .C(n14508), .D(n14507), 
        .Z(n14537) );
  HS65_LL_NAND4ABX3 U15747 ( .A(n14514), .B(n14513), .C(n14512), .D(n14511), 
        .Z(n14518) );
  HS65_LL_NOR3X1 U15748 ( .A(n14516), .B(n15317), .C(n14515), .Z(n14517) );
  HS65_LL_NAND4ABX3 U15749 ( .A(n14519), .B(n14518), .C(n14517), .D(n15278), 
        .Z(n14536) );
  HS65_LL_OAI112X1 U15750 ( .A(n14522), .B(n14521), .C(n14520), .D(n15299), 
        .Z(n14525) );
  HS65_LL_NAND4ABX3 U15751 ( .A(n14526), .B(n14525), .C(n14524), .D(n14523), 
        .Z(n14535) );
  HS65_LL_NOR4ABX2 U15752 ( .A(n14530), .B(n14529), .C(n14528), .D(n14527), 
        .Z(n14531) );
  HS65_LL_NAND3AX3 U15753 ( .A(n14533), .B(n14532), .C(n14531), .Z(n14534) );
  HS65_LL_MX41X4 U15754 ( .D0(n14537), .S0(n15328), .D1(n14536), .S1(n15326), 
        .D2(n14535), .S2(n15324), .D3(n14534), .S3(n15322), .Z(n15619) );
  HS65_LLS_XOR3X2 U15755 ( .A(n15277), .B(n15641), .C(n15619), .Z(n14538) );
  HS65_LL_MUX21I1X3 U15756 ( .D0(w2[31]), .D1(w2[31]), .S0(n14538), .Z(n14539)
         );
  HS65_LL_MUXI21X2 U15757 ( .D0(n15602), .D1(n15603), .S0(n14539), .Z(n14540)
         );
  HS65_LL_CBI4I1X3 U15758 ( .A(text_in_r[63]), .B(w2[31]), .C(n14541), .D(
        n14540), .Z(N153) );
  HS65_LL_IVX2 U15759 ( .A(n15113), .Z(n14552) );
  HS65_LL_MUXI21X2 U15760 ( .D0(n14552), .D1(n15113), .S0(n15531), .Z(n14643)
         );
  HS65_LLS_XOR3X2 U15761 ( .A(n15523), .B(n15347), .C(n14643), .Z(n14542) );
  HS65_LL_MUXI21X2 U15762 ( .D0(n14542), .D1(text_in_r[118]), .S0(n15545), .Z(
        n14543) );
  HS65_LLS_XNOR2X3 U15763 ( .A(w0[22]), .B(n14543), .Z(N264) );
  HS65_LL_MUXI21X2 U15764 ( .D0(n15123), .D1(n15124), .S0(n14544), .Z(n14545)
         );
  HS65_LL_MUXI21X2 U15765 ( .D0(n14857), .D1(n14858), .S0(n14545), .Z(n14546)
         );
  HS65_LL_OAI21X2 U15766 ( .A(n11557), .B(text_in_r[87]), .C(n14546), .Z(
        n14547) );
  HS65_LLS_XNOR2X3 U15767 ( .A(w1[23]), .B(n14547), .Z(N201) );
  HS65_LL_MUXI21X2 U15768 ( .D0(n15275), .D1(n15276), .S0(n14965), .Z(n14548)
         );
  HS65_LL_MUXI21X2 U15769 ( .D0(n14857), .D1(n14858), .S0(n14548), .Z(n14549)
         );
  HS65_LL_OAI21X2 U15770 ( .A(n11557), .B(text_in_r[72]), .C(n14549), .Z(
        n14550) );
  HS65_LLS_XNOR2X3 U15771 ( .A(w1[8]), .B(n14550), .Z(N178) );
  HS65_LL_OAI21X2 U15772 ( .A(w0[31]), .B(text_in_r[127]), .C(n14822), .Z(
        n14556) );
  HS65_LL_IVX2 U15773 ( .A(n15254), .Z(n15253) );
  HS65_LL_MUX21I1X3 U15774 ( .D0(w0[31]), .D1(w0[31]), .S0(n15253), .Z(n14551)
         );
  HS65_LL_MUXI21X2 U15775 ( .D0(n14552), .D1(n15113), .S0(n14551), .Z(n14553)
         );
  HS65_LL_MUXI21X2 U15776 ( .D0(n15251), .D1(n15252), .S0(n14553), .Z(n14554)
         );
  HS65_LL_MUXI21X2 U15777 ( .D0(n14798), .D1(n14797), .S0(n14554), .Z(n14555)
         );
  HS65_LL_CBI4I1X3 U15778 ( .A(text_in_r[127]), .B(w0[31]), .C(n14556), .D(
        n14555), .Z(N281) );
  HS65_LL_MUXI21X2 U15779 ( .D0(n15262), .D1(n15261), .S0(n14793), .Z(n14557)
         );
  HS65_LL_MUXI21X2 U15780 ( .D0(n14803), .D1(n14804), .S0(n14557), .Z(n14558)
         );
  HS65_LL_OAI21X2 U15781 ( .A(n11557), .B(text_in_r[120]), .C(n14558), .Z(
        n14559) );
  HS65_LLS_XNOR2X3 U15782 ( .A(w0[24]), .B(n14559), .Z(N274) );
  HS65_LL_OAI21X2 U15783 ( .A(w1[9]), .B(text_in_r[73]), .C(n15698), .Z(n14564) );
  HS65_LL_IVX2 U15784 ( .A(n15371), .Z(n15372) );
  HS65_LL_MUXI21X2 U15785 ( .D0(n15454), .D1(n15453), .S0(w1[9]), .Z(n14560)
         );
  HS65_LLS_XOR3X2 U15786 ( .A(n14961), .B(n15273), .C(n14560), .Z(n14561) );
  HS65_LL_MUXI21X2 U15787 ( .D0(n15371), .D1(n15372), .S0(n14561), .Z(n14562)
         );
  HS65_LL_MUXI21X2 U15788 ( .D0(n14858), .D1(n14857), .S0(n14562), .Z(n14563)
         );
  HS65_LL_CBI4I1X3 U15789 ( .A(text_in_r[73]), .B(w1[9]), .C(n14564), .D(
        n14563), .Z(N179) );
  HS65_LL_OAI21X2 U15790 ( .A(w3[25]), .B(text_in_r[25]), .C(n15734), .Z(
        n14620) );
  HS65_LL_NAND2X2 U15791 ( .A(n15214), .B(n14565), .Z(n14600) );
  HS65_LL_NOR4ABX2 U15792 ( .A(n14568), .B(n14567), .C(n14600), .D(n14566), 
        .Z(n14569) );
  HS65_LL_NAND3X2 U15793 ( .A(n14570), .B(n14587), .C(n14569), .Z(n14615) );
  HS65_LL_NAND4ABX3 U15794 ( .A(n14573), .B(n14572), .C(n14915), .D(n14571), 
        .Z(n14588) );
  HS65_LL_NOR2X2 U15795 ( .A(n14574), .B(n14595), .Z(n14576) );
  HS65_LL_NAND4ABX3 U15796 ( .A(n14923), .B(n14576), .C(n14575), .D(n15228), 
        .Z(n14578) );
  HS65_LL_NAND4ABX3 U15797 ( .A(n14579), .B(n14578), .C(n14577), .D(n14601), 
        .Z(n15198) );
  HS65_LL_NAND3X2 U15798 ( .A(n14582), .B(n14581), .C(n14580), .Z(n14583) );
  HS65_LL_AOI112X2 U15799 ( .A(n14585), .B(n14584), .C(n15198), .D(n14583), 
        .Z(n14586) );
  HS65_LL_NAND4ABX3 U15800 ( .A(n14589), .B(n14588), .C(n14587), .D(n14586), 
        .Z(n14614) );
  HS65_LL_NOR2X2 U15801 ( .A(n14591), .B(n14590), .Z(n14910) );
  HS65_LL_IVX2 U15802 ( .A(n14592), .Z(n15224) );
  HS65_LL_NOR2X2 U15803 ( .A(n15224), .B(n14593), .Z(n14605) );
  HS65_LL_NOR2X2 U15804 ( .A(n14595), .B(n14594), .Z(n14597) );
  HS65_LL_NOR4ABX2 U15805 ( .A(n14605), .B(n14598), .C(n14597), .D(n14596), 
        .Z(n14599) );
  HS65_LL_NAND4ABX3 U15806 ( .A(n14600), .B(n15232), .C(n14910), .D(n14599), 
        .Z(n14613) );
  HS65_LL_NAND4ABX3 U15807 ( .A(n14602), .B(n15209), .C(n15217), .D(n14601), 
        .Z(n14603) );
  HS65_LL_NOR4ABX2 U15808 ( .A(n15203), .B(n14605), .C(n14604), .D(n14603), 
        .Z(n14919) );
  HS65_LL_NOR4ABX2 U15809 ( .A(n14919), .B(n14607), .C(n15227), .D(n14606), 
        .Z(n14608) );
  HS65_LL_NAND4ABX3 U15810 ( .A(n14611), .B(n14610), .C(n14609), .D(n14608), 
        .Z(n14612) );
  HS65_LL_MX41X4 U15811 ( .D0(n14615), .S0(n15240), .D1(n14614), .S1(n15238), 
        .D2(n14613), .S2(n15236), .D3(n14612), .S3(n15234), .Z(n15714) );
  HS65_LLS_XNOR2X3 U15812 ( .A(n15343), .B(n15432), .Z(n15673) );
  HS65_LL_MUXI21X2 U15813 ( .D0(n15250), .D1(w3[25]), .S0(n15519), .Z(n14616)
         );
  HS65_LLS_XOR3X2 U15814 ( .A(n15673), .B(n15693), .C(n14616), .Z(n14617) );
  HS65_LL_MUX21I1X3 U15815 ( .D0(n15714), .D1(n15714), .S0(n14617), .Z(n14618)
         );
  HS65_LL_MUXI21X2 U15816 ( .D0(n15742), .D1(n15743), .S0(n14618), .Z(n14619)
         );
  HS65_LL_CBI4I1X3 U15817 ( .A(text_in_r[25]), .B(w3[25]), .C(n14620), .D(
        n14619), .Z(N83) );
  HS65_LL_OAI21X2 U15818 ( .A(w0[11]), .B(text_in_r[107]), .C(n14822), .Z(
        n14626) );
  HS65_LL_MUXI21X2 U15819 ( .D0(n15352), .D1(w0[11]), .S0(n15256), .Z(n14621)
         );
  HS65_LLS_XOR3X2 U15820 ( .A(n14819), .B(n14622), .C(n14621), .Z(n14623) );
  HS65_LL_MUXI21X2 U15821 ( .D0(n15353), .D1(n15354), .S0(n14623), .Z(n14624)
         );
  HS65_LL_MUXI21X2 U15822 ( .D0(n14798), .D1(n14797), .S0(n14624), .Z(n14625)
         );
  HS65_LL_CBI4I1X3 U15823 ( .A(text_in_r[107]), .B(w0[11]), .C(n14626), .D(
        n14625), .Z(N245) );
  HS65_LL_OAI21X2 U15824 ( .A(w2[27]), .B(text_in_r[59]), .C(n15688), .Z(
        n14632) );
  HS65_LLS_XOR3X2 U15825 ( .A(w2[27]), .B(n15607), .C(n14627), .Z(n14629) );
  HS65_LLS_XOR3X2 U15826 ( .A(n14629), .B(n15629), .C(n14628), .Z(n14630) );
  HS65_LL_MUXI21X2 U15827 ( .D0(n15651), .D1(n15652), .S0(n14630), .Z(n14631)
         );
  HS65_LL_CBI4I1X3 U15828 ( .A(text_in_r[59]), .B(w2[27]), .C(n14632), .D(
        n14631), .Z(N149) );
  HS65_LLS_XNOR2X3 U15829 ( .A(n15553), .B(n15261), .Z(n14788) );
  HS65_LLS_XOR3X2 U15830 ( .A(n15556), .B(n14633), .C(n14788), .Z(n14634) );
  HS65_LL_MUXI21X2 U15831 ( .D0(n14634), .D1(text_in_r[96]), .S0(n15545), .Z(
        n14635) );
  HS65_LLS_XNOR2X3 U15832 ( .A(w0[0]), .B(n14635), .Z(N226) );
  HS65_LL_OAI21X2 U15833 ( .A(w3[11]), .B(text_in_r[11]), .C(n14822), .Z(
        n14642) );
  HS65_LLS_XOR2X3 U15834 ( .A(n15740), .B(n15513), .Z(n14636) );
  HS65_LL_NOR2AX3 U15835 ( .A(n14636), .B(n15698), .Z(n15696) );
  HS65_LL_NOR2X2 U15836 ( .A(n14822), .B(n14636), .Z(n15695) );
  HS65_LL_IVX2 U15837 ( .A(n14815), .Z(n15340) );
  HS65_LLS_XOR3X2 U15838 ( .A(n15340), .B(n14638), .C(n14637), .Z(n14639) );
  HS65_LL_MUXI21X2 U15839 ( .D0(n15431), .D1(w3[11]), .S0(n14639), .Z(n14640)
         );
  HS65_LL_MUXI21X2 U15840 ( .D0(n15696), .D1(n15695), .S0(n14640), .Z(n14641)
         );
  HS65_LL_CBI4I1X3 U15841 ( .A(text_in_r[11]), .B(w3[11]), .C(n14642), .D(
        n14641), .Z(N53) );
  HS65_LL_IVX2 U15842 ( .A(n15345), .Z(n15346) );
  HS65_LL_MUXI21X2 U15843 ( .D0(n15346), .D1(n15345), .S0(n14643), .Z(n14644)
         );
  HS65_LL_MUXI21X2 U15844 ( .D0(n14803), .D1(n14804), .S0(n14644), .Z(n14645)
         );
  HS65_LL_OAI21X2 U15845 ( .A(n11557), .B(text_in_r[103]), .C(n14645), .Z(
        n14646) );
  HS65_LLS_XNOR2X3 U15846 ( .A(w0[7]), .B(n14646), .Z(N233) );
  HS65_LL_OAI21X2 U15847 ( .A(w1[27]), .B(text_in_r[91]), .C(n15727), .Z(
        n14698) );
  HS65_LL_IVX2 U15848 ( .A(w1[27]), .Z(n15132) );
  HS65_LLS_XNOR2X3 U15849 ( .A(n14647), .B(n15133), .Z(n14960) );
  HS65_LL_NOR4ABX2 U15850 ( .A(n14651), .B(n14650), .C(n14649), .D(n14648), 
        .Z(n14653) );
  HS65_LL_NAND4ABX3 U15851 ( .A(n14655), .B(n14654), .C(n14653), .D(n14652), 
        .Z(n14692) );
  HS65_LL_AOI112X2 U15852 ( .A(n14659), .B(n14658), .C(n14657), .D(n14656), 
        .Z(n14662) );
  HS65_LL_NOR4ABX2 U15853 ( .A(n14663), .B(n14662), .C(n14661), .D(n14660), 
        .Z(n14688) );
  HS65_LL_NOR4ABX2 U15854 ( .A(n14667), .B(n14666), .C(n14665), .D(n14664), 
        .Z(n14672) );
  HS65_LL_NOR3X1 U15855 ( .A(n14670), .B(n14669), .C(n14668), .Z(n14671) );
  HS65_LL_NAND3X2 U15856 ( .A(n14673), .B(n14672), .C(n14671), .Z(n14684) );
  HS65_LL_NOR4ABX2 U15857 ( .A(n14677), .B(n14676), .C(n14675), .D(n14674), 
        .Z(n14678) );
  HS65_LL_NAND4ABX3 U15858 ( .A(n14681), .B(n14680), .C(n14679), .D(n14678), 
        .Z(n14682) );
  HS65_LL_AOI22X1 U15859 ( .A(n14685), .B(n14684), .C(n14683), .D(n14682), .Z(
        n14686) );
  HS65_LL_CBI4I1X3 U15860 ( .A(n14689), .B(n14688), .C(n14687), .D(n14686), 
        .Z(n14690) );
  HS65_LL_CBI4I6X2 U15861 ( .A(n14693), .B(n14692), .C(n14691), .D(n14690), 
        .Z(n15449) );
  HS65_LLS_XOR3X2 U15862 ( .A(n14960), .B(n15449), .C(n14694), .Z(n14695) );
  HS65_LL_MUXI21X2 U15863 ( .D0(n15132), .D1(w1[27]), .S0(n14695), .Z(n14696)
         );
  HS65_LL_MUXI21X2 U15864 ( .D0(n14843), .D1(n14842), .S0(n14696), .Z(n14697)
         );
  HS65_LL_CBI4I1X3 U15865 ( .A(text_in_r[91]), .B(w1[27]), .C(n14698), .D(
        n14697), .Z(N213) );
  HS65_LL_OAI21X2 U15866 ( .A(w3[9]), .B(text_in_r[9]), .C(n14822), .Z(n14754)
         );
  HS65_LL_NOR4ABX2 U15867 ( .A(n14702), .B(n14701), .C(n14700), .D(n14699), 
        .Z(n14704) );
  HS65_LL_NAND4ABX3 U15868 ( .A(n14706), .B(n14705), .C(n14704), .D(n14703), 
        .Z(n14749) );
  HS65_LL_NOR4ABX2 U15869 ( .A(n14710), .B(n14709), .C(n14708), .D(n14707), 
        .Z(n14715) );
  HS65_LL_NOR4ABX2 U15870 ( .A(n14713), .B(n14728), .C(n14712), .D(n14711), 
        .Z(n14714) );
  HS65_LL_NAND4ABX3 U15871 ( .A(n14717), .B(n14716), .C(n14715), .D(n14714), 
        .Z(n14747) );
  HS65_LL_NOR3X1 U15872 ( .A(n14719), .B(n14740), .C(n14718), .Z(n14721) );
  HS65_LL_OAI112X1 U15873 ( .A(n14723), .B(n14722), .C(n14721), .D(n14720), 
        .Z(n14726) );
  HS65_LL_NAND4ABX3 U15874 ( .A(n14727), .B(n14726), .C(n14725), .D(n14724), 
        .Z(n14745) );
  HS65_LL_NAND2X2 U15875 ( .A(n14729), .B(n14728), .Z(n14730) );
  HS65_LL_AOI112X2 U15876 ( .A(n14733), .B(n14732), .C(n14731), .D(n14730), 
        .Z(n14739) );
  HS65_LL_NOR4ABX2 U15877 ( .A(n14737), .B(n14736), .C(n14735), .D(n14734), 
        .Z(n14738) );
  HS65_LL_NAND4ABX3 U15878 ( .A(n14741), .B(n14740), .C(n14739), .D(n14738), 
        .Z(n14743) );
  HS65_LL_MX41X4 U15879 ( .D0(n14749), .S0(n14748), .D1(n14747), .S1(n14746), 
        .D2(n14745), .S2(n14744), .D3(n14743), .S3(n14742), .Z(n15656) );
  HS65_LL_IVX2 U15880 ( .A(n15656), .Z(n15657) );
  HS65_LLS_XOR3X2 U15881 ( .A(n15343), .B(w3[9]), .C(n15719), .Z(n14750) );
  HS65_LL_MUXI21X2 U15882 ( .D0(n15667), .D1(n15434), .S0(n14750), .Z(n14751)
         );
  HS65_LL_MUXI21X2 U15883 ( .D0(n15656), .D1(n15657), .S0(n14751), .Z(n14752)
         );
  HS65_LL_MUXI21X2 U15884 ( .D0(n15696), .D1(n15695), .S0(n14752), .Z(n14753)
         );
  HS65_LL_CBI4I1X3 U15885 ( .A(text_in_r[9]), .B(w3[9]), .C(n14754), .D(n14753), .Z(N51) );
  HS65_LL_OAI21X2 U15886 ( .A(w1[12]), .B(text_in_r[76]), .C(n15727), .Z(
        n14759) );
  HS65_LL_IVX2 U15887 ( .A(w1[12]), .Z(n15364) );
  HS65_LL_MUXI21X2 U15888 ( .D0(w1[12]), .D1(n15364), .S0(n15449), .Z(n14755)
         );
  HS65_LLS_XOR3X2 U15889 ( .A(n14952), .B(n15269), .C(n14755), .Z(n14756) );
  HS65_LL_MUX21I1X3 U15890 ( .D0(n15365), .D1(n15365), .S0(n14756), .Z(n14757)
         );
  HS65_LL_MUXI21X2 U15891 ( .D0(n14858), .D1(n14857), .S0(n14757), .Z(n14758)
         );
  HS65_LL_CBI4I1X3 U15892 ( .A(text_in_r[76]), .B(w1[12]), .C(n14759), .D(
        n14758), .Z(N182) );
  HS65_LL_OAI21X2 U15893 ( .A(w3[27]), .B(text_in_r[27]), .C(n15727), .Z(
        n14765) );
  HS65_LLS_XNOR2X3 U15894 ( .A(n15247), .B(n15342), .Z(n15718) );
  HS65_LLS_XOR3X2 U15895 ( .A(n14761), .B(n14760), .C(n15718), .Z(n14762) );
  HS65_LL_MUXI21X2 U15896 ( .D0(n15246), .D1(w3[27]), .S0(n14762), .Z(n14763)
         );
  HS65_LL_MUXI21X2 U15897 ( .D0(n15742), .D1(n15743), .S0(n14763), .Z(n14764)
         );
  HS65_LL_CBI4I1X3 U15898 ( .A(text_in_r[27]), .B(w3[27]), .C(n14765), .D(
        n14764), .Z(N85) );
  HS65_LLS_XNOR2X3 U15899 ( .A(n15254), .B(n15347), .Z(n14979) );
  HS65_LL_MUXI21X2 U15900 ( .D0(n15111), .D1(n15112), .S0(n14979), .Z(n14766)
         );
  HS65_LL_MUXI21X2 U15901 ( .D0(n14797), .D1(n14798), .S0(n14766), .Z(n14767)
         );
  HS65_LL_OAI21X2 U15902 ( .A(n11557), .B(text_in_r[119]), .C(n14767), .Z(
        n14768) );
  HS65_LLS_XNOR2X3 U15903 ( .A(w0[23]), .B(n14768), .Z(N265) );
  HS65_LL_OAI21X2 U15904 ( .A(w0[27]), .B(text_in_r[123]), .C(n14822), .Z(
        n14773) );
  HS65_LLS_XOR3X2 U15905 ( .A(w0[27]), .B(n14831), .C(n14769), .Z(n14770) );
  HS65_LLS_XOR3X2 U15906 ( .A(n15119), .B(n15258), .C(n14770), .Z(n14771) );
  HS65_LL_MUXI21X2 U15907 ( .D0(n14804), .D1(n14803), .S0(n14771), .Z(n14772)
         );
  HS65_LL_CBI4I1X3 U15908 ( .A(text_in_r[123]), .B(w0[27]), .C(n14773), .D(
        n14772), .Z(N277) );
  HS65_LLS_XOR2X3 U15909 ( .A(n14788), .B(n15551), .Z(n14774) );
  HS65_LL_MUXI21X2 U15910 ( .D0(n14797), .D1(n14798), .S0(n14774), .Z(n14775)
         );
  HS65_LL_OAI21X2 U15911 ( .A(n11557), .B(text_in_r[104]), .C(n14775), .Z(
        n14776) );
  HS65_LLS_XNOR2X3 U15912 ( .A(w0[8]), .B(n14776), .Z(N242) );
  HS65_LL_MUX21I1X3 U15913 ( .D0(n15131), .D1(n15131), .S0(n15449), .Z(n14853)
         );
  HS65_LL_IVX2 U15914 ( .A(w1[19]), .Z(n15272) );
  HS65_LL_MUXI21X2 U15915 ( .D0(n15272), .D1(w1[19]), .S0(n15365), .Z(n14777)
         );
  HS65_LLS_XOR3X2 U15916 ( .A(n14853), .B(n14778), .C(n14777), .Z(n14782) );
  HS65_LL_OAI21X2 U15917 ( .A(n14964), .B(n14782), .C(n14832), .Z(n14781) );
  HS65_LL_IVX2 U15918 ( .A(text_in_r[83]), .Z(n14779) );
  HS65_LL_OAI212X3 U15919 ( .A(w1[19]), .B(text_in_r[83]), .C(n15272), .D(
        n14779), .E(n15545), .Z(n14780) );
  HS65_LL_CBI4I1X3 U15920 ( .A(n14782), .B(n14964), .C(n14781), .D(n14780), 
        .Z(N197) );
  HS65_LL_IVX2 U15921 ( .A(w1[4]), .Z(n15448) );
  HS65_LL_MUXI21X2 U15922 ( .D0(n15448), .D1(w1[4]), .S0(n15129), .Z(n14783)
         );
  HS65_LLS_XOR3X2 U15923 ( .A(n14853), .B(n14973), .C(n14783), .Z(n14787) );
  HS65_LLS_XNOR2X3 U15924 ( .A(n15363), .B(n15269), .Z(n14985) );
  HS65_LL_OAI21X2 U15925 ( .A(n14985), .B(n14787), .C(n14832), .Z(n14786) );
  HS65_LL_IVX2 U15926 ( .A(text_in_r[68]), .Z(n14784) );
  HS65_LL_OAI212X3 U15927 ( .A(w1[4]), .B(text_in_r[68]), .C(n15448), .D(
        n14784), .E(n15698), .Z(n14785) );
  HS65_LL_CBI4I1X3 U15928 ( .A(n14787), .B(n14985), .C(n14786), .D(n14785), 
        .Z(N166) );
  HS65_LL_OAI21X2 U15929 ( .A(w0[25]), .B(text_in_r[121]), .C(n14822), .Z(
        n14792) );
  HS65_LL_IVX2 U15930 ( .A(w0[25]), .Z(n15121) );
  HS65_LLS_XOR2X3 U15931 ( .A(n15259), .B(n15355), .Z(n15557) );
  HS65_LLS_XOR3X2 U15932 ( .A(n15557), .B(n14788), .C(n15441), .Z(n14789) );
  HS65_LL_MUXI21X2 U15933 ( .D0(n15121), .D1(w0[25]), .S0(n14789), .Z(n14790)
         );
  HS65_LL_MUXI21X2 U15934 ( .D0(n14804), .D1(n14803), .S0(n14790), .Z(n14791)
         );
  HS65_LL_CBI4I1X3 U15935 ( .A(text_in_r[121]), .B(w0[25]), .C(n14792), .D(
        n14791), .Z(N275) );
  HS65_LL_OAI21X2 U15936 ( .A(w0[9]), .B(text_in_r[105]), .C(n15727), .Z(
        n14800) );
  HS65_LLS_XOR3X2 U15937 ( .A(n14794), .B(n15259), .C(n14793), .Z(n14795) );
  HS65_LL_MUXI21X2 U15938 ( .D0(n15356), .D1(w0[9]), .S0(n14795), .Z(n14796)
         );
  HS65_LL_MUXI21X2 U15939 ( .D0(n14798), .D1(n14797), .S0(n14796), .Z(n14799)
         );
  HS65_LL_CBI4I1X3 U15940 ( .A(text_in_r[105]), .B(w0[9]), .C(n14800), .D(
        n14799), .Z(N243) );
  HS65_LL_OAI21X2 U15941 ( .A(w0[28]), .B(text_in_r[124]), .C(n14822), .Z(
        n14806) );
  HS65_LLS_XOR3X2 U15942 ( .A(w0[28]), .B(n14976), .C(n15540), .Z(n14801) );
  HS65_LLS_XOR3X2 U15943 ( .A(n15256), .B(n15117), .C(n14801), .Z(n14802) );
  HS65_LL_MUXI21X2 U15944 ( .D0(n14804), .D1(n14803), .S0(n14802), .Z(n14805)
         );
  HS65_LL_CBI4I1X3 U15945 ( .A(text_in_r[124]), .B(w0[28]), .C(n14806), .D(
        n14805), .Z(N278) );
  HS65_LLS_XOR2X3 U15946 ( .A(n15714), .B(n15656), .Z(n15692) );
  HS65_LL_IVX2 U15947 ( .A(w3[1]), .Z(n15520) );
  HS65_LL_MUXI21X2 U15948 ( .D0(n15520), .D1(w3[1]), .S0(n15249), .Z(n14807)
         );
  HS65_LLS_XOR3X2 U15949 ( .A(n15692), .B(n14807), .C(n15713), .Z(n14812) );
  HS65_LL_OAI21X2 U15950 ( .A(n15673), .B(n14812), .C(n14808), .Z(n14811) );
  HS65_LL_IVX2 U15951 ( .A(text_in_r[1]), .Z(n14809) );
  HS65_LL_OAI212X3 U15952 ( .A(w3[1]), .B(text_in_r[1]), .C(n15520), .D(n14809), .E(n15698), .Z(n14810) );
  HS65_LL_CBI4I1X3 U15953 ( .A(n14812), .B(n15673), .C(n14811), .D(n14810), 
        .Z(N35) );
  HS65_LL_OAI21X2 U15954 ( .A(w3[28]), .B(text_in_r[28]), .C(n15734), .Z(
        n14818) );
  HS65_LL_MUXI21X2 U15955 ( .D0(w3[28]), .D1(n15244), .S0(n15514), .Z(n14813)
         );
  HS65_LLS_XOR3X2 U15956 ( .A(n15678), .B(n15245), .C(n14813), .Z(n14814) );
  HS65_LL_MUXI21X2 U15957 ( .D0(n14815), .D1(n15340), .S0(n14814), .Z(n14816)
         );
  HS65_LL_MUXI21X2 U15958 ( .D0(n15742), .D1(n15743), .S0(n14816), .Z(n14817)
         );
  HS65_LL_CBI4I1X3 U15959 ( .A(text_in_r[28]), .B(w3[28]), .C(n14818), .D(
        n14817), .Z(N86) );
  HS65_LLS_XNOR2X3 U15960 ( .A(n15119), .B(n14819), .Z(n15535) );
  HS65_LLS_XOR3X2 U15961 ( .A(n15354), .B(n15557), .C(n15535), .Z(n14820) );
  HS65_LL_MUXI21X2 U15962 ( .D0(n14820), .D1(text_in_r[114]), .S0(n15545), .Z(
        n14821) );
  HS65_LLS_XNOR2X3 U15963 ( .A(w0[18]), .B(n14821), .Z(N260) );
  HS65_LL_OAI21X2 U15964 ( .A(w3[12]), .B(text_in_r[12]), .C(n14822), .Z(
        n14829) );
  HS65_LL_IVX2 U15965 ( .A(n14826), .Z(n15430) );
  HS65_LL_MUXI21X2 U15966 ( .D0(n14823), .D1(n15514), .S0(n15243), .Z(n15725)
         );
  HS65_LL_MUXI21X2 U15967 ( .D0(n15429), .D1(w3[12]), .S0(n15516), .Z(n14824)
         );
  HS65_LLS_XOR3X2 U15968 ( .A(n15338), .B(n15725), .C(n14824), .Z(n14825) );
  HS65_LL_MUXI21X2 U15969 ( .D0(n14826), .D1(n15430), .S0(n14825), .Z(n14827)
         );
  HS65_LL_MUXI21X2 U15970 ( .D0(n15696), .D1(n15695), .S0(n14827), .Z(n14828)
         );
  HS65_LL_CBI4I1X3 U15971 ( .A(text_in_r[12]), .B(w3[12]), .C(n14829), .D(
        n14828), .Z(N54) );
  HS65_LL_MUXI21X2 U15972 ( .D0(w0[3]), .D1(n15440), .S0(n15117), .Z(n14830)
         );
  HS65_LLS_XOR3X2 U15973 ( .A(n14831), .B(n14830), .C(n15535), .Z(n14836) );
  HS65_LL_OAI21X2 U15974 ( .A(n15556), .B(n14836), .C(n14832), .Z(n14835) );
  HS65_LL_IVX2 U15975 ( .A(text_in_r[99]), .Z(n14833) );
  HS65_LL_OAI212X3 U15976 ( .A(w0[3]), .B(text_in_r[99]), .C(n15440), .D(
        n14833), .E(n15545), .Z(n14834) );
  HS65_LL_CBI4I1X3 U15977 ( .A(n14836), .B(n15556), .C(n14835), .D(n14834), 
        .Z(N229) );
  HS65_LL_OAI21X2 U15978 ( .A(w1[28]), .B(text_in_r[92]), .C(n15698), .Z(
        n14845) );
  HS65_LL_IVX2 U15979 ( .A(n15271), .Z(n14840) );
  HS65_LL_IVX2 U15980 ( .A(w1[28]), .Z(n15130) );
  HS65_LL_MUXI21X2 U15981 ( .D0(n15130), .D1(w1[28]), .S0(n14837), .Z(n14838)
         );
  HS65_LLS_XOR3X2 U15982 ( .A(n14985), .B(n15131), .C(n14838), .Z(n14839) );
  HS65_LL_MUXI21X2 U15983 ( .D0(n14840), .D1(n15271), .S0(n14839), .Z(n14841)
         );
  HS65_LL_MUXI21X2 U15984 ( .D0(n14843), .D1(n14842), .S0(n14841), .Z(n14844)
         );
  HS65_LL_CBI4I1X3 U15985 ( .A(text_in_r[92]), .B(w1[28]), .C(n14845), .D(
        n14844), .Z(N214) );
  HS65_LL_OAI21X2 U15986 ( .A(w2[11]), .B(text_in_r[43]), .C(n15688), .Z(
        n14851) );
  HS65_LL_IVX2 U15987 ( .A(w2[11]), .Z(n15422) );
  HS65_LL_MUXI21X2 U15988 ( .D0(w2[11]), .D1(n15422), .S0(n15510), .Z(n14846)
         );
  HS65_LLS_XOR3X2 U15989 ( .A(n14847), .B(n15331), .C(n14846), .Z(n14848) );
  HS65_LL_MUXI21X2 U15990 ( .D0(n15423), .D1(n15424), .S0(n14848), .Z(n14849)
         );
  HS65_LL_MUXI21X2 U15991 ( .D0(n15602), .D1(n15603), .S0(n14849), .Z(n14850)
         );
  HS65_LL_CBI4I1X3 U15992 ( .A(text_in_r[43]), .B(w2[11]), .C(n14851), .D(
        n14850), .Z(N117) );
  HS65_LL_OAI21X2 U15993 ( .A(w1[11]), .B(text_in_r[75]), .C(n15698), .Z(
        n14860) );
  HS65_LL_IVX2 U15994 ( .A(w1[11]), .Z(n15366) );
  HS65_LL_MUXI21X2 U15995 ( .D0(n15366), .D1(w1[11]), .S0(n15271), .Z(n14852)
         );
  HS65_LLS_XOR3X2 U15996 ( .A(n14854), .B(n14853), .C(n14852), .Z(n14855) );
  HS65_LL_MUXI21X2 U15997 ( .D0(n15367), .D1(n15368), .S0(n14855), .Z(n14856)
         );
  HS65_LL_MUXI21X2 U15998 ( .D0(n14858), .D1(n14857), .S0(n14856), .Z(n14859)
         );
  HS65_LL_CBI4I1X3 U15999 ( .A(text_in_r[75]), .B(w1[11]), .C(n14860), .D(
        n14859), .Z(N181) );
  HS65_LL_OAI21X2 U16000 ( .A(w3[31]), .B(text_in_r[31]), .C(n15734), .Z(
        n14945) );
  HS65_LL_NAND3X2 U16001 ( .A(n14862), .B(n14861), .C(n14886), .Z(n14869) );
  HS65_LL_NOR4ABX2 U16002 ( .A(n14866), .B(n14865), .C(n14864), .D(n14863), 
        .Z(n14868) );
  HS65_LL_NAND4ABX3 U16003 ( .A(n14870), .B(n14869), .C(n14868), .D(n14867), 
        .Z(n14900) );
  HS65_LL_NOR4ABX2 U16004 ( .A(n14874), .B(n14873), .C(n14872), .D(n14871), 
        .Z(n14897) );
  HS65_LL_NOR3X1 U16005 ( .A(n14877), .B(n14876), .C(n14875), .Z(n14896) );
  HS65_LL_NOR4ABX2 U16006 ( .A(n14881), .B(n14880), .C(n14879), .D(n14878), 
        .Z(n14882) );
  HS65_LL_NAND4ABX3 U16007 ( .A(n14885), .B(n14884), .C(n14883), .D(n14882), 
        .Z(n14892) );
  HS65_LL_NAND4ABX3 U16008 ( .A(n14889), .B(n14888), .C(n14887), .D(n14886), 
        .Z(n14890) );
  HS65_LL_AOI22X1 U16009 ( .A(n14893), .B(n14892), .C(n14891), .D(n14890), .Z(
        n14894) );
  HS65_LL_CBI4I1X3 U16010 ( .A(n14897), .B(n14896), .C(n14895), .D(n14894), 
        .Z(n14898) );
  HS65_LL_CBI4I6X2 U16011 ( .A(n14901), .B(n14900), .C(n14899), .D(n14898), 
        .Z(n15662) );
  HS65_LL_IVX2 U16012 ( .A(n15662), .Z(n15708) );
  HS65_LL_NOR4ABX2 U16013 ( .A(n14937), .B(n14904), .C(n14903), .D(n14902), 
        .Z(n14906) );
  HS65_LL_NAND4ABX3 U16014 ( .A(n14908), .B(n14907), .C(n14906), .D(n14905), 
        .Z(n14939) );
  HS65_LL_NAND3X2 U16015 ( .A(n14911), .B(n14910), .C(n14909), .Z(n14912) );
  HS65_LL_NOR4ABX2 U16016 ( .A(n14915), .B(n14914), .C(n14913), .D(n14912), 
        .Z(n14936) );
  HS65_LL_NOR3AX2 U16017 ( .A(n14918), .B(n14917), .C(n14916), .Z(n15201) );
  HS65_LL_NAND4ABX3 U16018 ( .A(n14921), .B(n14920), .C(n14919), .D(n15201), 
        .Z(n14933) );
  HS65_LL_NOR2X2 U16019 ( .A(n14923), .B(n14922), .Z(n15220) );
  HS65_LL_CBI4I6X2 U16020 ( .A(sa03[7]), .B(n14925), .C(n14924), .D(sa03[6]), 
        .Z(n14926) );
  HS65_LL_NOR4ABX2 U16021 ( .A(n14929), .B(n14928), .C(n14927), .D(n14926), 
        .Z(n14930) );
  HS65_LL_NAND3X2 U16022 ( .A(n14931), .B(n15220), .C(n14930), .Z(n14932) );
  HS65_LL_AOI22X1 U16023 ( .A(n15240), .B(n14933), .C(n15236), .D(n14932), .Z(
        n14934) );
  HS65_LL_CBI4I1X3 U16024 ( .A(n14937), .B(n14936), .C(n14935), .D(n14934), 
        .Z(n14938) );
  HS65_LL_CBI4I6X2 U16025 ( .A(n14940), .B(n14939), .C(n15234), .D(n14938), 
        .Z(n15733) );
  HS65_LL_MUXI21X2 U16026 ( .D0(n15708), .D1(n15662), .S0(n15733), .Z(n14941)
         );
  HS65_LL_MUX21I1X3 U16027 ( .D0(n15337), .D1(n15337), .S0(n14941), .Z(n14942)
         );
  HS65_LL_MUXI21X2 U16028 ( .D0(n15195), .D1(w3[31]), .S0(n14942), .Z(n14943)
         );
  HS65_LL_MUXI21X2 U16029 ( .D0(n15696), .D1(n15695), .S0(n14943), .Z(n14944)
         );
  HS65_LL_CBI4I1X3 U16030 ( .A(text_in_r[31]), .B(w3[31]), .C(n14945), .D(
        n14944), .Z(N89) );
  HS65_LLS_XOR3X2 U16031 ( .A(n15609), .B(n14946), .C(n15423), .Z(n14947) );
  HS65_LL_MUXI21X2 U16032 ( .D0(n14947), .D1(text_in_r[50]), .S0(n15734), .Z(
        n14948) );
  HS65_LLS_XNOR2X3 U16033 ( .A(w2[18]), .B(n14948), .Z(N132) );
  HS65_LLS_XOR3X2 U16034 ( .A(n14984), .B(n15359), .C(n14949), .Z(n14950) );
  HS65_LL_MUXI21X2 U16035 ( .D0(n14950), .D1(text_in_r[70]), .S0(n15688), .Z(
        n14951) );
  HS65_LLS_XNOR2X3 U16036 ( .A(w1[6]), .B(n14951), .Z(N168) );
  HS65_LLS_XOR3X2 U16037 ( .A(n14952), .B(n14956), .C(n15127), .Z(n14953) );
  HS65_LL_MUXI21X2 U16038 ( .D0(n14953), .D1(text_in_r[69]), .S0(n15688), .Z(
        n14954) );
  HS65_LLS_XNOR2X3 U16039 ( .A(w1[5]), .B(n14954), .Z(N167) );
  HS65_LLS_XOR3X2 U16040 ( .A(n14957), .B(n14956), .C(n14955), .Z(n14958) );
  HS65_LL_MUXI21X2 U16041 ( .D0(n14958), .D1(text_in_r[86]), .S0(n15688), .Z(
        n14959) );
  HS65_LLS_XNOR2X3 U16042 ( .A(w1[22]), .B(n14959), .Z(N200) );
  HS65_LLS_XOR3X2 U16043 ( .A(n14961), .B(n14960), .C(n15367), .Z(n14962) );
  HS65_LL_MUXI21X2 U16044 ( .D0(n14962), .D1(text_in_r[66]), .S0(n15688), .Z(
        n14963) );
  HS65_LLS_XNOR2X3 U16045 ( .A(w1[2]), .B(n14963), .Z(N164) );
  HS65_LLS_XOR3X2 U16046 ( .A(n14965), .B(n14964), .C(n15371), .Z(n14966) );
  HS65_LL_MUXI21X2 U16047 ( .D0(n14966), .D1(text_in_r[80]), .S0(n15688), .Z(
        n14967) );
  HS65_LLS_XNOR2X3 U16048 ( .A(w1[16]), .B(n14967), .Z(N194) );
  HS65_LLS_XOR3X2 U16049 ( .A(n14969), .B(n14968), .C(n15367), .Z(n14970) );
  HS65_LL_MUXI21X2 U16050 ( .D0(n14970), .D1(text_in_r[82]), .S0(n15688), .Z(
        n14971) );
  HS65_LLS_XNOR2X3 U16051 ( .A(w1[18]), .B(n14971), .Z(N196) );
  HS65_LLS_XOR3X2 U16052 ( .A(n14973), .B(n14972), .C(n15137), .Z(n14974) );
  HS65_LL_MUXI21X2 U16053 ( .D0(n14974), .D1(text_in_r[64]), .S0(n15688), .Z(
        n14975) );
  HS65_LLS_XNOR2X3 U16054 ( .A(w1[0]), .B(n14975), .Z(N162) );
  HS65_LL_IVX2 U16055 ( .A(n15115), .Z(n15114) );
  HS65_LL_MUXI21X2 U16056 ( .D0(n15114), .D1(n15115), .S0(n15521), .Z(n15542)
         );
  HS65_LLS_XOR3X2 U16057 ( .A(n15349), .B(n14976), .C(n15542), .Z(n14977) );
  HS65_LL_MUXI21X2 U16058 ( .D0(n14977), .D1(text_in_r[117]), .S0(n15688), .Z(
        n14978) );
  HS65_LLS_XNOR2X3 U16059 ( .A(w0[21]), .B(n14978), .Z(N263) );
  HS65_LL_MUXI21X2 U16060 ( .D0(n15114), .D1(n15115), .S0(n14979), .Z(n15529)
         );
  HS65_LLS_XNOR2X3 U16061 ( .A(n15529), .B(n14980), .Z(n14981) );
  HS65_LL_MUXI21X2 U16062 ( .D0(n14981), .D1(text_in_r[102]), .S0(n15688), .Z(
        n14982) );
  HS65_LLS_XNOR2X3 U16063 ( .A(w0[6]), .B(n14982), .Z(N232) );
  HS65_LLS_XOR3X2 U16064 ( .A(n14985), .B(n14984), .C(n14983), .Z(n14986) );
  HS65_LL_MUXI21X2 U16065 ( .D0(n14986), .D1(text_in_r[85]), .S0(n15688), .Z(
        n14987) );
  HS65_LLS_XNOR2X3 U16066 ( .A(w1[21]), .B(n14987), .Z(N199) );
  HS65_LL_NOR2AX3 U16067 ( .A(n14989), .B(n14988), .Z(n15748) );
  HS65_LL_NAND3X2 U16068 ( .A(n14990), .B(n15748), .C(n14996), .Z(n15004) );
  HS65_LL_NAND4ABX3 U16069 ( .A(\u0/r0/rcnt [0]), .B(\u0/r0/rcnt [1]), .C(
        \u0/r0/N81 ), .D(n14992), .Z(n14997) );
  HS65_LL_OAI21X2 U16070 ( .A(n14991), .B(n15004), .C(n14997), .Z(\u0/r0/N75 )
         );
  HS65_LL_NOR2X2 U16071 ( .A(\u0/r0/rcnt [3]), .B(n14996), .Z(n14993) );
  HS65_LL_NAND3X2 U16072 ( .A(\u0/r0/rcnt [0]), .B(n14993), .C(n15844), .Z(
        n15747) );
  HS65_LL_OAI21X2 U16073 ( .A(n15748), .B(n15747), .C(n14997), .Z(\u0/r0/N72 )
         );
  HS65_LL_NAND2X2 U16074 ( .A(\u0/r0/N78 ), .B(n14992), .Z(n15000) );
  HS65_LL_IVX2 U16075 ( .A(n14993), .Z(n14995) );
  HS65_LL_NAND2X2 U16076 ( .A(n14999), .B(n15108), .Z(n14994) );
  HS65_LL_OAI21X2 U16077 ( .A(n15000), .B(n14995), .C(n14994), .Z(\u0/r0/N73 )
         );
  HS65_LL_IVX2 U16078 ( .A(n14996), .Z(n15001) );
  HS65_LL_IVX2 U16079 ( .A(n14997), .Z(n14998) );
  HS65_LL_AOI12X2 U16080 ( .A(n14999), .B(n15844), .C(n14998), .Z(n15002) );
  HS65_LL_OAI21X2 U16081 ( .A(n15001), .B(n15000), .C(n15002), .Z(\u0/r0/N71 )
         );
  HS65_LL_NAND2X2 U16082 ( .A(\u0/r0/rcnt [0]), .B(n15844), .Z(n15003) );
  HS65_LL_OAI21X2 U16083 ( .A(n15004), .B(n15003), .C(n15002), .Z(\u0/r0/N74 )
         );
  HS65_LLS_XNOR2X3 U16084 ( .A(w1[21]), .B(n15005), .Z(n15830) );
  HS65_LL_OAI21X2 U16085 ( .A(w2[21]), .B(n15830), .C(n15108), .Z(n15006) );
  HS65_LL_AOI12X2 U16086 ( .A(w2[21]), .B(n15830), .C(n15006), .Z(n15790) );
  HS65_LL_AO12X4 U16087 ( .A(n15110), .B(key[53]), .C(n15790), .Z(\u0/N195 )
         );
  HS65_LLS_XNOR2X3 U16088 ( .A(w1[23]), .B(n15007), .Z(n15832) );
  HS65_LL_OAI21X2 U16089 ( .A(w2[23]), .B(n15832), .C(n15108), .Z(n15008) );
  HS65_LL_AOI12X2 U16090 ( .A(w2[23]), .B(n15832), .C(n15008), .Z(n15794) );
  HS65_LL_AO12X4 U16091 ( .A(n15110), .B(key[55]), .C(n15794), .Z(\u0/N197 )
         );
  HS65_LL_IVX4 U16092 ( .A(n15806), .Z(n15826) );
  HS65_LL_MUXI21X2 U16093 ( .D0(w1[11]), .D1(n15366), .S0(n15009), .Z(n15820)
         );
  HS65_LL_OAI21X2 U16094 ( .A(w2[11]), .B(n15820), .C(n15843), .Z(n15010) );
  HS65_LL_AOI12X2 U16095 ( .A(w2[11]), .B(n15820), .C(n15010), .Z(n15771) );
  HS65_LL_AO12X4 U16096 ( .A(n15826), .B(key[43]), .C(n15771), .Z(\u0/N185 )
         );
  HS65_LL_MUXI21X2 U16097 ( .D0(w1[20]), .D1(n15270), .S0(n15011), .Z(n15829)
         );
  HS65_LL_OAI21X2 U16098 ( .A(w2[20]), .B(n15829), .C(n15108), .Z(n15012) );
  HS65_LL_AOI12X2 U16099 ( .A(w2[20]), .B(n15829), .C(n15012), .Z(n15788) );
  HS65_LL_AO12X4 U16100 ( .A(n15110), .B(key[52]), .C(n15788), .Z(\u0/N194 )
         );
  HS65_LL_MUXI21X2 U16101 ( .D0(w1[15]), .D1(n15014), .S0(n15013), .Z(n15823)
         );
  HS65_LL_OAI21X2 U16102 ( .A(w2[15]), .B(n15823), .C(n15843), .Z(n15015) );
  HS65_LL_AOI12X2 U16103 ( .A(w2[15]), .B(n15823), .C(n15015), .Z(n15777) );
  HS65_LL_AO12X4 U16104 ( .A(n15826), .B(key[47]), .C(n15777), .Z(\u0/N189 )
         );
  HS65_LLS_XNOR2X3 U16105 ( .A(n15016), .B(w1[5]), .Z(n15814) );
  HS65_LL_OAI21X2 U16106 ( .A(w2[5]), .B(n15814), .C(n15108), .Z(n15017) );
  HS65_LL_AOI12X2 U16107 ( .A(w2[5]), .B(n15814), .C(n15017), .Z(n15759) );
  HS65_LL_AO12X4 U16108 ( .A(n15842), .B(key[37]), .C(n15759), .Z(\u0/N179 )
         );
  HS65_LL_MUXI21X2 U16109 ( .D0(w1[12]), .D1(n15364), .S0(n15018), .Z(n15821)
         );
  HS65_LL_OAI21X2 U16110 ( .A(w2[12]), .B(n15821), .C(n15843), .Z(n15019) );
  HS65_LL_AOI12X2 U16111 ( .A(w2[12]), .B(n15821), .C(n15019), .Z(n15773) );
  HS65_LL_AO12X4 U16112 ( .A(n15826), .B(key[44]), .C(n15773), .Z(\u0/N186 )
         );
  HS65_LL_MUXI21X2 U16113 ( .D0(w1[17]), .D1(n15274), .S0(n15020), .Z(n15825)
         );
  HS65_LL_OAI21X2 U16114 ( .A(w2[17]), .B(n15825), .C(n15843), .Z(n15021) );
  HS65_LL_AOI12X2 U16115 ( .A(w2[17]), .B(n15825), .C(n15021), .Z(n15781) );
  HS65_LL_AO12X4 U16116 ( .A(n15110), .B(key[49]), .C(n15781), .Z(\u0/N191 )
         );
  HS65_LL_MUXI21X2 U16117 ( .D0(w1[14]), .D1(n15360), .S0(n15022), .Z(n15822)
         );
  HS65_LL_OAI21X2 U16118 ( .A(w2[14]), .B(n15822), .C(n15843), .Z(n15023) );
  HS65_LL_AOI12X2 U16119 ( .A(w2[14]), .B(n15822), .C(n15023), .Z(n15775) );
  HS65_LL_AO12X4 U16120 ( .A(n15826), .B(key[46]), .C(n15775), .Z(\u0/N188 )
         );
  HS65_LLS_XNOR2X3 U16121 ( .A(w1[2]), .B(n15024), .Z(n15811) );
  HS65_LL_OAI21X2 U16122 ( .A(w2[2]), .B(n15811), .C(n15844), .Z(n15025) );
  HS65_LL_AOI12X2 U16123 ( .A(w2[2]), .B(n15811), .C(n15025), .Z(n15753) );
  HS65_LL_AO12X4 U16124 ( .A(n15842), .B(key[34]), .C(n15753), .Z(\u0/N176 )
         );
  HS65_LLS_XNOR2X3 U16125 ( .A(n15026), .B(w1[8]), .Z(n15817) );
  HS65_LL_OAI21X2 U16126 ( .A(w2[8]), .B(n15817), .C(n15843), .Z(n15027) );
  HS65_LL_AOI12X2 U16127 ( .A(w2[8]), .B(n15817), .C(n15027), .Z(n15765) );
  HS65_LL_AO12X4 U16128 ( .A(n15842), .B(key[40]), .C(n15765), .Z(\u0/N182 )
         );
  HS65_LLS_XNOR2X3 U16129 ( .A(n15028), .B(w1[22]), .Z(n15831) );
  HS65_LL_OAI21X2 U16130 ( .A(w2[22]), .B(n15831), .C(n15108), .Z(n15029) );
  HS65_LL_AOI12X2 U16131 ( .A(w2[22]), .B(n15831), .C(n15029), .Z(n15792) );
  HS65_LL_AO12X4 U16132 ( .A(n15110), .B(key[54]), .C(n15792), .Z(\u0/N196 )
         );
  HS65_LL_IVX2 U16133 ( .A(w1[9]), .Z(n15370) );
  HS65_LL_MUXI21X2 U16134 ( .D0(w1[9]), .D1(n15370), .S0(n15030), .Z(n15818)
         );
  HS65_LL_OAI21X2 U16135 ( .A(w2[9]), .B(n15818), .C(n15843), .Z(n15031) );
  HS65_LL_AOI12X2 U16136 ( .A(w2[9]), .B(n15818), .C(n15031), .Z(n15767) );
  HS65_LL_AO12X4 U16137 ( .A(n15842), .B(key[41]), .C(n15767), .Z(\u0/N183 )
         );
  HS65_LL_MUXI21X2 U16138 ( .D0(w1[1]), .D1(n15452), .S0(n15032), .Z(n15810)
         );
  HS65_LL_OAI21X2 U16139 ( .A(w2[1]), .B(n15810), .C(n15108), .Z(n15033) );
  HS65_LL_AOI12X2 U16140 ( .A(w2[1]), .B(n15810), .C(n15033), .Z(n15751) );
  HS65_LL_AO12X4 U16141 ( .A(n15842), .B(key[33]), .C(n15751), .Z(\u0/N175 )
         );
  HS65_LL_MUXI21X2 U16142 ( .D0(w1[10]), .D1(n15035), .S0(n15034), .Z(n15819)
         );
  HS65_LL_OAI21X2 U16143 ( .A(w2[10]), .B(n15819), .C(n15843), .Z(n15036) );
  HS65_LL_AOI12X2 U16144 ( .A(w2[10]), .B(n15819), .C(n15036), .Z(n15769) );
  HS65_LL_AO12X4 U16145 ( .A(n15842), .B(key[42]), .C(n15769), .Z(\u0/N184 )
         );
  HS65_LL_MUXI21X2 U16146 ( .D0(w1[19]), .D1(n15272), .S0(n15037), .Z(n15828)
         );
  HS65_LL_OAI21X2 U16147 ( .A(w2[19]), .B(n15828), .C(n15108), .Z(n15038) );
  HS65_LL_AOI12X2 U16148 ( .A(w2[19]), .B(n15828), .C(n15038), .Z(n15786) );
  HS65_LL_AO12X4 U16149 ( .A(n15110), .B(key[51]), .C(n15786), .Z(\u0/N193 )
         );
  HS65_LLS_XNOR2X3 U16150 ( .A(n15039), .B(w1[7]), .Z(n15816) );
  HS65_LL_OAI21X2 U16151 ( .A(w2[7]), .B(n15816), .C(n15843), .Z(n15040) );
  HS65_LL_AOI12X2 U16152 ( .A(w2[7]), .B(n15816), .C(n15040), .Z(n15763) );
  HS65_LL_AO12X4 U16153 ( .A(n15842), .B(key[39]), .C(n15763), .Z(\u0/N181 )
         );
  HS65_LLS_XNOR2X3 U16154 ( .A(n15041), .B(w1[0]), .Z(n15809) );
  HS65_LL_OAI21X2 U16155 ( .A(w2[0]), .B(n15809), .C(n15108), .Z(n15042) );
  HS65_LL_AOI12X2 U16156 ( .A(w2[0]), .B(n15809), .C(n15042), .Z(n15749) );
  HS65_LL_AO12X4 U16157 ( .A(n15842), .B(key[32]), .C(n15749), .Z(\u0/N174 )
         );
  HS65_LL_MUXI21X2 U16158 ( .D0(w1[4]), .D1(n15448), .S0(n15043), .Z(n15813)
         );
  HS65_LL_OAI21X2 U16159 ( .A(w2[4]), .B(n15813), .C(n15108), .Z(n15044) );
  HS65_LL_AOI12X2 U16160 ( .A(w2[4]), .B(n15813), .C(n15044), .Z(n15757) );
  HS65_LL_AO12X4 U16161 ( .A(n15826), .B(key[36]), .C(n15757), .Z(\u0/N178 )
         );
  HS65_LL_CBI4I1X3 U16162 ( .A(n15048), .B(n15047), .C(n15046), .D(n15045), 
        .Z(n15055) );
  HS65_LL_NOR4ABX2 U16163 ( .A(n15052), .B(n15051), .C(n15050), .D(n15049), 
        .Z(n15053) );
  HS65_LL_NAND4ABX3 U16164 ( .A(n15056), .B(n15055), .C(n15054), .D(n15053), 
        .Z(n15089) );
  HS65_LL_NOR2X2 U16165 ( .A(n15058), .B(n15057), .Z(n15059) );
  HS65_LL_NAND4ABX3 U16166 ( .A(n15062), .B(n15061), .C(n15060), .D(n15059), 
        .Z(n15065) );
  HS65_LL_NAND4ABX3 U16167 ( .A(n15066), .B(n15065), .C(n15064), .D(n15063), 
        .Z(n15087) );
  HS65_LL_NOR4ABX2 U16168 ( .A(n15070), .B(n15069), .C(n15068), .D(n15067), 
        .Z(n15071) );
  HS65_LL_NAND4ABX3 U16169 ( .A(n15073), .B(n15076), .C(n15072), .D(n15071), 
        .Z(n15085) );
  HS65_LL_NAND4ABX3 U16170 ( .A(n15077), .B(n15076), .C(n15075), .D(n15074), 
        .Z(n15080) );
  HS65_LL_NAND4ABX3 U16171 ( .A(n15081), .B(n15080), .C(n15079), .D(n15078), 
        .Z(n15083) );
  HS65_LL_MX41X4 U16172 ( .D0(n15089), .S0(n15088), .D1(n15087), .S1(n15086), 
        .D2(n15085), .S2(n15084), .D3(n15083), .S3(n15082), .Z(n15090) );
  HS65_LLS_XOR3X2 U16173 ( .A(\u0/rcon [31]), .B(w0[31]), .C(n15090), .Z(
        n15840) );
  HS65_LL_MUXI21X2 U16174 ( .D0(n15091), .D1(w1[31]), .S0(n15840), .Z(n15838)
         );
  HS65_LL_OAI21X2 U16175 ( .A(w2[31]), .B(n15838), .C(n15108), .Z(n15092) );
  HS65_LL_AOI12X2 U16176 ( .A(w2[31]), .B(n15838), .C(n15092), .Z(n15807) );
  HS65_LL_AO12X4 U16177 ( .A(n15842), .B(key[63]), .C(n15807), .Z(\u0/N205 )
         );
  HS65_LL_MUXI21X2 U16178 ( .D0(w1[3]), .D1(n15450), .S0(n15093), .Z(n15812)
         );
  HS65_LL_OAI21X2 U16179 ( .A(w2[3]), .B(n15812), .C(n15108), .Z(n15094) );
  HS65_LL_AOI12X2 U16180 ( .A(w2[3]), .B(n15812), .C(n15094), .Z(n15755) );
  HS65_LL_AO12X4 U16181 ( .A(n15842), .B(key[35]), .C(n15755), .Z(\u0/N177 )
         );
  HS65_LLS_XNOR2X3 U16182 ( .A(w1[16]), .B(n15095), .Z(n15824) );
  HS65_LL_OAI21X2 U16183 ( .A(w2[16]), .B(n15824), .C(n15843), .Z(n15096) );
  HS65_LL_AOI12X2 U16184 ( .A(w2[16]), .B(n15824), .C(n15096), .Z(n15779) );
  HS65_LL_AO12X4 U16185 ( .A(n15842), .B(key[48]), .C(n15779), .Z(\u0/N190 )
         );
  HS65_LLS_XNOR2X3 U16186 ( .A(n15097), .B(w1[6]), .Z(n15815) );
  HS65_LL_OAI21X2 U16187 ( .A(w2[6]), .B(n15815), .C(n15108), .Z(n15098) );
  HS65_LL_AOI12X2 U16188 ( .A(w2[6]), .B(n15815), .C(n15098), .Z(n15761) );
  HS65_LL_AO12X4 U16189 ( .A(n15842), .B(key[38]), .C(n15761), .Z(\u0/N180 )
         );
  HS65_LL_MUXI21X2 U16190 ( .D0(w1[28]), .D1(n15130), .S0(n15099), .Z(n15836)
         );
  HS65_LL_OAI21X2 U16191 ( .A(w2[28]), .B(n15836), .C(n15108), .Z(n15100) );
  HS65_LL_AOI12X2 U16192 ( .A(w2[28]), .B(n15836), .C(n15100), .Z(n15802) );
  HS65_LL_AO12X4 U16193 ( .A(n15783), .B(key[60]), .C(n15802), .Z(\u0/N202 )
         );
  HS65_LL_MUXI21X2 U16194 ( .D0(w1[30]), .D1(n15126), .S0(n15101), .Z(n15837)
         );
  HS65_LL_OAI21X2 U16195 ( .A(w2[30]), .B(n15837), .C(n15108), .Z(n15102) );
  HS65_LL_AOI12X2 U16196 ( .A(w2[30]), .B(n15837), .C(n15102), .Z(n15804) );
  HS65_LL_AO12X4 U16197 ( .A(n15842), .B(key[62]), .C(n15804), .Z(\u0/N204 )
         );
  HS65_LLS_XNOR2X3 U16198 ( .A(n15103), .B(w1[24]), .Z(n15833) );
  HS65_LL_OAI21X2 U16199 ( .A(w2[24]), .B(n15833), .C(n15108), .Z(n15104) );
  HS65_LL_AOI12X2 U16200 ( .A(w2[24]), .B(n15833), .C(n15104), .Z(n15796) );
  HS65_LL_AO12X4 U16201 ( .A(n15110), .B(key[56]), .C(n15796), .Z(\u0/N198 )
         );
  HS65_LL_MUXI21X2 U16202 ( .D0(w1[27]), .D1(n15132), .S0(n15105), .Z(n15835)
         );
  HS65_LL_OAI21X2 U16203 ( .A(w2[27]), .B(n15835), .C(n15108), .Z(n15106) );
  HS65_LL_AOI12X2 U16204 ( .A(w2[27]), .B(n15835), .C(n15106), .Z(n15800) );
  HS65_LL_AO12X4 U16205 ( .A(n15783), .B(key[59]), .C(n15800), .Z(\u0/N201 )
         );
  HS65_LL_MUXI21X2 U16206 ( .D0(w1[26]), .D1(n15134), .S0(n15107), .Z(n15834)
         );
  HS65_LL_OAI21X2 U16207 ( .A(w2[26]), .B(n15834), .C(n15108), .Z(n15109) );
  HS65_LL_AOI12X2 U16208 ( .A(w2[26]), .B(n15834), .C(n15109), .Z(n15798) );
  HS65_LL_AO12X4 U16209 ( .A(n15110), .B(key[58]), .C(n15798), .Z(\u0/N200 )
         );
  HS65_LL_MUXI21X2 U16210 ( .D0(n15112), .D1(n15111), .S0(w0[31]), .Z(N378) );
  HS65_LL_IVX2 U16211 ( .A(w0[30]), .Z(n15534) );
  HS65_LL_MUXI21X2 U16212 ( .D0(w0[30]), .D1(n15534), .S0(n15113), .Z(N379) );
  HS65_LL_MUXI21X2 U16213 ( .D0(n15115), .D1(n15114), .S0(w0[29]), .Z(N380) );
  HS65_LL_IVX2 U16214 ( .A(w0[28]), .Z(n15116) );
  HS65_LL_MUXI21X2 U16215 ( .D0(n15116), .D1(w0[28]), .S0(n15524), .Z(N381) );
  HS65_LL_IVX2 U16216 ( .A(w0[27]), .Z(n15118) );
  HS65_LL_MUXI21X2 U16217 ( .D0(n15118), .D1(w0[27]), .S0(n15117), .Z(N382) );
  HS65_LL_MUXI21X2 U16218 ( .D0(w0[26]), .D1(n15120), .S0(n15119), .Z(N383) );
  HS65_LL_MUXI21X2 U16219 ( .D0(n15121), .D1(w0[25]), .S0(n15552), .Z(N384) );
  HS65_LL_IVX2 U16220 ( .A(n15553), .Z(n15122) );
  HS65_LL_MUXI21X2 U16221 ( .D0(n15122), .D1(n15553), .S0(w0[24]), .Z(N385) );
  HS65_LL_MUXI21X2 U16222 ( .D0(n15124), .D1(n15123), .S0(w1[31]), .Z(N386) );
  HS65_LL_MUXI21X2 U16223 ( .D0(w1[30]), .D1(n15126), .S0(n15125), .Z(N387) );
  HS65_LL_MUXI21X2 U16224 ( .D0(n15128), .D1(w1[29]), .S0(n15127), .Z(N388) );
  HS65_LL_MUXI21X2 U16225 ( .D0(n15130), .D1(w1[28]), .S0(n15129), .Z(N389) );
  HS65_LL_MUXI21X2 U16226 ( .D0(n15132), .D1(w1[27]), .S0(n15131), .Z(N390) );
  HS65_LL_MUXI21X2 U16227 ( .D0(n15134), .D1(w1[26]), .S0(n15133), .Z(N391) );
  HS65_LL_MUXI21X2 U16228 ( .D0(n15136), .D1(w1[25]), .S0(n15135), .Z(N392) );
  HS65_LL_IVX2 U16229 ( .A(n15137), .Z(n15138) );
  HS65_LL_MUXI21X2 U16230 ( .D0(n15138), .D1(n15137), .S0(w1[24]), .Z(N393) );
  HS65_LL_MUXI21X2 U16231 ( .D0(n15593), .D1(n15594), .S0(w2[31]), .Z(N394) );
  HS65_LL_IVX2 U16232 ( .A(w2[30]), .Z(n15577) );
  HS65_LL_MUXI21X2 U16233 ( .D0(n15577), .D1(w2[30]), .S0(n15641), .Z(N395) );
  HS65_LL_NAND3X2 U16234 ( .A(n15141), .B(n15140), .C(n15139), .Z(n15142) );
  HS65_LL_NOR4ABX2 U16235 ( .A(n15145), .B(n15144), .C(n15143), .D(n15142), 
        .Z(n15146) );
  HS65_LL_NAND3X2 U16236 ( .A(n15148), .B(n15147), .C(n15146), .Z(n15187) );
  HS65_LL_NOR4ABX2 U16237 ( .A(n15151), .B(n15150), .C(n15171), .D(n15149), 
        .Z(n15157) );
  HS65_LL_NOR4ABX2 U16238 ( .A(n15155), .B(n15154), .C(n15153), .D(n15152), 
        .Z(n15156) );
  HS65_LL_NAND4ABX3 U16239 ( .A(n15159), .B(n15158), .C(n15157), .D(n15156), 
        .Z(n15185) );
  HS65_LL_NOR4ABX2 U16240 ( .A(n15163), .B(n15162), .C(n15161), .D(n15160), 
        .Z(n15164) );
  HS65_LL_NAND4ABX3 U16241 ( .A(n15167), .B(n15166), .C(n15165), .D(n15164), 
        .Z(n15183) );
  HS65_LL_NAND4ABX3 U16242 ( .A(n15171), .B(n15170), .C(n15169), .D(n15168), 
        .Z(n15179) );
  HS65_LL_NAND4ABX3 U16243 ( .A(n15175), .B(n15174), .C(n15173), .D(n15172), 
        .Z(n15178) );
  HS65_LL_NAND4ABX3 U16244 ( .A(n15179), .B(n15178), .C(n15177), .D(n15176), 
        .Z(n15181) );
  HS65_LL_MX41X4 U16245 ( .D0(n15187), .S0(n15186), .D1(n15185), .S1(n15184), 
        .D2(n15183), .S2(n15182), .D3(n15181), .S3(n15180), .Z(n15614) );
  HS65_LL_IVX2 U16246 ( .A(n15614), .Z(n15613) );
  HS65_LL_MUXI21X2 U16247 ( .D0(n15613), .D1(n15614), .S0(w2[29]), .Z(N396) );
  HS65_LL_IVX2 U16248 ( .A(w2[28]), .Z(n15188) );
  HS65_LL_MUXI21X2 U16249 ( .D0(n15188), .D1(w2[28]), .S0(n15568), .Z(N397) );
  HS65_LL_IVX2 U16250 ( .A(w2[27]), .Z(n15190) );
  HS65_LL_MUXI21X2 U16251 ( .D0(n15190), .D1(w2[27]), .S0(n15189), .Z(N398) );
  HS65_LL_IVX2 U16252 ( .A(w2[26]), .Z(n15191) );
  HS65_LL_MUXI21X2 U16253 ( .D0(n15191), .D1(w2[26]), .S0(n15629), .Z(N399) );
  HS65_LL_MUXI21X2 U16254 ( .D0(n15193), .D1(w2[25]), .S0(n15192), .Z(N400) );
  HS65_LL_IVX2 U16255 ( .A(w2[24]), .Z(n15566) );
  HS65_LL_MUXI21X2 U16256 ( .D0(w2[24]), .D1(n15566), .S0(n15625), .Z(N401) );
  HS65_LL_MUXI21X2 U16257 ( .D0(n15195), .D1(w3[31]), .S0(n15194), .Z(N402) );
  HS65_LL_MUXI21X2 U16258 ( .D0(w3[30]), .D1(n15666), .S0(n15733), .Z(N403) );
  HS65_LL_NAND4ABX3 U16259 ( .A(n15225), .B(n15197), .C(n15217), .D(n15196), 
        .Z(n15204) );
  HS65_LL_NOR4ABX2 U16260 ( .A(n15201), .B(n15200), .C(n15199), .D(n15198), 
        .Z(n15202) );
  HS65_LL_NAND4ABX3 U16261 ( .A(n15205), .B(n15204), .C(n15203), .D(n15202), 
        .Z(n15241) );
  HS65_LL_NAND4ABX3 U16262 ( .A(n15209), .B(n15208), .C(n15207), .D(n15206), 
        .Z(n15210) );
  HS65_LL_NOR3X1 U16263 ( .A(n15211), .B(n15223), .C(n15210), .Z(n15212) );
  HS65_LL_NAND3X2 U16264 ( .A(n15214), .B(n15213), .C(n15212), .Z(n15239) );
  HS65_LL_NOR4ABX2 U16265 ( .A(n15218), .B(n15217), .C(n15216), .D(n15215), 
        .Z(n15219) );
  HS65_LL_NAND4ABX3 U16266 ( .A(n15222), .B(n15221), .C(n15220), .D(n15219), 
        .Z(n15237) );
  HS65_LL_NOR3X1 U16267 ( .A(n15225), .B(n15224), .C(n15223), .Z(n15231) );
  HS65_LL_NOR4ABX2 U16268 ( .A(n15229), .B(n15228), .C(n15227), .D(n15226), 
        .Z(n15230) );
  HS65_LL_NAND4ABX3 U16269 ( .A(n15233), .B(n15232), .C(n15231), .D(n15230), 
        .Z(n15235) );
  HS65_LL_MX41X4 U16270 ( .D0(n15241), .S0(n15240), .D1(n15239), .S1(n15238), 
        .D2(n15237), .S2(n15236), .D3(n15235), .S3(n15234), .Z(n15703) );
  HS65_LL_IVX2 U16271 ( .A(n15703), .Z(n15702) );
  HS65_LL_MUXI21X2 U16272 ( .D0(w3[29]), .D1(n15242), .S0(n15702), .Z(N404) );
  HS65_LL_MUXI21X2 U16273 ( .D0(w3[28]), .D1(n15244), .S0(n15243), .Z(N405) );
  HS65_LL_MUXI21X2 U16274 ( .D0(n15246), .D1(w3[27]), .S0(n15245), .Z(N406) );
  HS65_LL_MUXI21X2 U16275 ( .D0(n15248), .D1(w3[26]), .S0(n15247), .Z(N407) );
  HS65_LL_MUXI21X2 U16276 ( .D0(w3[25]), .D1(n15250), .S0(n15249), .Z(N408) );
  HS65_LL_MUXI21X2 U16277 ( .D0(n15661), .D1(w3[24]), .S0(n15714), .Z(N409) );
  HS65_LL_MUXI21X2 U16278 ( .D0(n15252), .D1(n15251), .S0(w0[23]), .Z(N410) );
  HS65_LL_MUXI21X2 U16279 ( .D0(n15254), .D1(n15253), .S0(w0[22]), .Z(N411) );
  HS65_LL_IVX2 U16280 ( .A(n15549), .Z(n15548) );
  HS65_LL_MUXI21X2 U16281 ( .D0(n15548), .D1(n15549), .S0(w0[21]), .Z(N412) );
  HS65_LL_MUXI21X2 U16282 ( .D0(n15255), .D1(w0[20]), .S0(n15522), .Z(N413) );
  HS65_LL_MUXI21X2 U16283 ( .D0(w0[19]), .D1(n15257), .S0(n15256), .Z(N414) );
  HS65_LL_IVX2 U16284 ( .A(n15258), .Z(n15537) );
  HS65_LL_MUXI21X2 U16285 ( .D0(n15537), .D1(n15258), .S0(w0[18]), .Z(N415) );
  HS65_LL_MUXI21X2 U16286 ( .D0(n15260), .D1(w0[17]), .S0(n15259), .Z(N416) );
  HS65_LL_MUXI21X2 U16287 ( .D0(n15262), .D1(n15261), .S0(w0[16]), .Z(N417) );
  HS65_LL_MUXI21X2 U16288 ( .D0(n15264), .D1(n15263), .S0(w1[23]), .Z(N418) );
  HS65_LL_MUXI21X2 U16289 ( .D0(n15266), .D1(n15265), .S0(w1[22]), .Z(N419) );
  HS65_LL_IVX2 U16290 ( .A(n15267), .Z(n15268) );
  HS65_LL_MUXI21X2 U16291 ( .D0(n15268), .D1(n15267), .S0(w1[21]), .Z(N420) );
  HS65_LL_MUXI21X2 U16292 ( .D0(n15270), .D1(w1[20]), .S0(n15269), .Z(N421) );
  HS65_LL_MUXI21X2 U16293 ( .D0(w1[19]), .D1(n15272), .S0(n15271), .Z(N422) );
  HS65_LL_MUXI21X2 U16294 ( .D0(n15274), .D1(w1[17]), .S0(n15273), .Z(N424) );
  HS65_LL_MUXI21X2 U16295 ( .D0(n15276), .D1(n15275), .S0(w1[16]), .Z(N425) );
  HS65_LL_IVX2 U16296 ( .A(w2[23]), .Z(n15598) );
  HS65_LL_MUXI21X2 U16297 ( .D0(n15598), .D1(w2[23]), .S0(n15277), .Z(N426) );
  HS65_LL_IVX2 U16298 ( .A(w2[22]), .Z(n15592) );
  HS65_LL_MUXI21X2 U16299 ( .D0(n15592), .D1(w2[22]), .S0(n15619), .Z(N427) );
  HS65_LL_IVX2 U16300 ( .A(w2[21]), .Z(n15586) );
  HS65_LL_NAND4ABX3 U16301 ( .A(n15280), .B(n15279), .C(n15278), .D(n15305), 
        .Z(n15284) );
  HS65_LL_OAI13X1 U16302 ( .A(sa13[1]), .B(n15282), .C(n15281), .D(n15319), 
        .Z(n15283) );
  HS65_LL_NOR3X1 U16303 ( .A(n15285), .B(n15284), .C(n15283), .Z(n15286) );
  HS65_LL_NAND3X2 U16304 ( .A(n15288), .B(n15287), .C(n15286), .Z(n15329) );
  HS65_LL_NOR4ABX2 U16305 ( .A(n15291), .B(n15290), .C(n15289), .D(n15317), 
        .Z(n15294) );
  HS65_LL_NOR4ABX2 U16306 ( .A(n15295), .B(n15294), .C(n15293), .D(n15292), 
        .Z(n15297) );
  HS65_LL_NAND3X2 U16307 ( .A(n15298), .B(n15297), .C(n15296), .Z(n15327) );
  HS65_LL_NAND3X2 U16308 ( .A(n15301), .B(n15300), .C(n15299), .Z(n15312) );
  HS65_LL_NOR4ABX2 U16309 ( .A(n15305), .B(n15304), .C(n15303), .D(n15302), 
        .Z(n15308) );
  HS65_LL_NOR4ABX2 U16310 ( .A(n15309), .B(n15308), .C(n15307), .D(n15306), 
        .Z(n15310) );
  HS65_LL_NAND4ABX3 U16311 ( .A(n15313), .B(n15312), .C(n15311), .D(n15310), 
        .Z(n15325) );
  HS65_LL_NAND4ABX3 U16312 ( .A(n15317), .B(n15316), .C(n15315), .D(n15314), 
        .Z(n15320) );
  HS65_LL_NAND4ABX3 U16313 ( .A(n15321), .B(n15320), .C(n15319), .D(n15318), 
        .Z(n15323) );
  HS65_LL_MX41X4 U16314 ( .D0(n15329), .S0(n15328), .D1(n15327), .S1(n15326), 
        .D2(n15325), .S2(n15324), .D3(n15323), .S3(n15322), .Z(n15575) );
  HS65_LL_IVX2 U16315 ( .A(n15575), .Z(n15616) );
  HS65_LL_MUXI21X2 U16316 ( .D0(w2[21]), .D1(n15586), .S0(n15616), .Z(N428) );
  HS65_LL_IVX2 U16317 ( .A(w2[20]), .Z(n15330) );
  HS65_LL_MUXI21X2 U16318 ( .D0(n15330), .D1(w2[20]), .S0(n15569), .Z(N429) );
  HS65_LL_MUXI21X2 U16319 ( .D0(n15332), .D1(w2[19]), .S0(n15331), .Z(N430) );
  HS65_LL_IVX2 U16320 ( .A(n15607), .Z(n15333) );
  HS65_LL_MUXI21X2 U16321 ( .D0(n15333), .D1(n15607), .S0(w2[18]), .Z(N431) );
  HS65_LL_MUXI21X2 U16322 ( .D0(n15335), .D1(n15334), .S0(w2[17]), .Z(N432) );
  HS65_LL_IVX2 U16323 ( .A(w2[16]), .Z(n15582) );
  HS65_LL_MUXI21X2 U16324 ( .D0(w2[16]), .D1(n15582), .S0(n15336), .Z(N433) );
  HS65_LL_MUXI21X2 U16325 ( .D0(n15691), .D1(w3[23]), .S0(n15337), .Z(N434) );
  HS65_LL_MUXI21X2 U16326 ( .D0(w3[22]), .D1(n15687), .S0(n15662), .Z(N435) );
  HS65_LL_IVX2 U16327 ( .A(n15664), .Z(n15705) );
  HS65_LL_MUXI21X2 U16328 ( .D0(w3[21]), .D1(n15681), .S0(n15705), .Z(N436) );
  HS65_LL_MUXI21X2 U16329 ( .D0(w3[20]), .D1(n15339), .S0(n15338), .Z(N437) );
  HS65_LL_MUXI21X2 U16330 ( .D0(w3[19]), .D1(n15341), .S0(n15340), .Z(N438) );
  HS65_LL_MUXI21X2 U16331 ( .D0(n15785), .D1(w3[18]), .S0(n15342), .Z(N439) );
  HS65_LL_MUXI21X2 U16332 ( .D0(w3[17]), .D1(n15344), .S0(n15343), .Z(N440) );
  HS65_LL_MUXI21X2 U16333 ( .D0(n15671), .D1(w3[16]), .S0(n15693), .Z(N441) );
  HS65_LL_MUXI21X2 U16334 ( .D0(n15346), .D1(n15345), .S0(w0[15]), .Z(N442) );
  HS65_LL_MUXI21X2 U16335 ( .D0(n15348), .D1(w0[14]), .S0(n15347), .Z(N443) );
  HS65_LL_MUXI21X2 U16336 ( .D0(w0[13]), .D1(n15541), .S0(n15349), .Z(N444) );
  HS65_LL_MUXI21X2 U16337 ( .D0(n15350), .D1(w0[12]), .S0(n15543), .Z(N445) );
  HS65_LL_MUXI21X2 U16338 ( .D0(n15352), .D1(w0[11]), .S0(n15351), .Z(N446) );
  HS65_LL_MUXI21X2 U16339 ( .D0(n15354), .D1(n15353), .S0(w0[10]), .Z(N447) );
  HS65_LL_MUXI21X2 U16340 ( .D0(n15356), .D1(w0[9]), .S0(n15355), .Z(N448) );
  HS65_LL_MUXI21X2 U16341 ( .D0(n15358), .D1(n15357), .S0(w1[15]), .Z(N450) );
  HS65_LL_MUXI21X2 U16342 ( .D0(w1[14]), .D1(n15360), .S0(n15359), .Z(N451) );
  HS65_LL_MUXI21X2 U16343 ( .D0(w1[13]), .D1(n15362), .S0(n15361), .Z(N452) );
  HS65_LL_MUXI21X2 U16344 ( .D0(w1[12]), .D1(n15364), .S0(n15363), .Z(N453) );
  HS65_LL_MUXI21X2 U16345 ( .D0(n15366), .D1(w1[11]), .S0(n15365), .Z(N454) );
  HS65_LL_MUXI21X2 U16346 ( .D0(n15368), .D1(n15367), .S0(w1[10]), .Z(N455) );
  HS65_LL_MUXI21X2 U16347 ( .D0(n15370), .D1(w1[9]), .S0(n15369), .Z(N456) );
  HS65_LL_MUXI21X2 U16348 ( .D0(n15372), .D1(n15371), .S0(w1[8]), .Z(N457) );
  HS65_LL_MUXI21X2 U16349 ( .D0(n15648), .D1(n15649), .S0(w2[15]), .Z(N458) );
  HS65_LL_IVX2 U16350 ( .A(w2[14]), .Z(n15622) );
  HS65_LL_MUXI21X2 U16351 ( .D0(w2[14]), .D1(n15622), .S0(n15574), .Z(N459) );
  HS65_LL_NAND4ABX3 U16352 ( .A(n15376), .B(n15375), .C(n15374), .D(n15373), 
        .Z(n15379) );
  HS65_LL_NAND4ABX3 U16353 ( .A(n15380), .B(n15379), .C(n15378), .D(n15377), 
        .Z(n15417) );
  HS65_LL_NAND4ABX3 U16354 ( .A(n15384), .B(n15383), .C(n15382), .D(n15381), 
        .Z(n15390) );
  HS65_LL_NAND4ABX3 U16355 ( .A(n15388), .B(n15387), .C(n15386), .D(n15385), 
        .Z(n15389) );
  HS65_LL_NOR4ABX2 U16356 ( .A(n15397), .B(n15391), .C(n15390), .D(n15389), 
        .Z(n15414) );
  HS65_LL_NAND4ABX3 U16357 ( .A(n15395), .B(n15394), .C(n15393), .D(n15392), 
        .Z(n15403) );
  HS65_LL_NAND4ABX3 U16358 ( .A(n15399), .B(n15398), .C(n15397), .D(n15396), 
        .Z(n15401) );
  HS65_LL_OAI13X1 U16359 ( .A(n15403), .B(n15402), .C(n15401), .D(n15400), .Z(
        n15412) );
  HS65_LL_NAND4ABX3 U16360 ( .A(n15407), .B(n15406), .C(n15405), .D(n15404), 
        .Z(n15409) );
  HS65_LL_OAI21X2 U16361 ( .A(n15410), .B(n15409), .C(n15408), .Z(n15411) );
  HS65_LL_OAI112X1 U16362 ( .A(n15414), .B(n15413), .C(n15412), .D(n15411), 
        .Z(n15415) );
  HS65_LL_CBI4I6X2 U16363 ( .A(n15418), .B(n15417), .C(n15416), .D(n15415), 
        .Z(n15637) );
  HS65_LL_IVX2 U16364 ( .A(n15637), .Z(n15567) );
  HS65_LL_MUXI21X2 U16365 ( .D0(n15637), .D1(n15567), .S0(w2[13]), .Z(N460) );
  HS65_LL_MUXI21X2 U16366 ( .D0(n15420), .D1(n15419), .S0(w2[12]), .Z(N461) );
  HS65_LL_MUXI21X2 U16367 ( .D0(n15422), .D1(w2[11]), .S0(n15421), .Z(N462) );
  HS65_LL_MUXI21X2 U16368 ( .D0(n15424), .D1(n15423), .S0(w2[10]), .Z(N463) );
  HS65_LL_MUXI21X2 U16369 ( .D0(n15426), .D1(n15425), .S0(w2[9]), .Z(N464) );
  HS65_LL_IVX2 U16370 ( .A(w2[8]), .Z(n15606) );
  HS65_LL_MUXI21X2 U16371 ( .D0(n15606), .D1(w2[8]), .S0(n15578), .Z(N465) );
  HS65_LL_MUXI21X2 U16372 ( .D0(w3[15]), .D1(n15427), .S0(n15739), .Z(N466) );
  HS65_LL_MUXI21X2 U16373 ( .D0(w3[14]), .D1(n15711), .S0(n15663), .Z(N467) );
  HS65_LL_MUXI21X2 U16374 ( .D0(w3[13]), .D1(n15707), .S0(n15726), .Z(N468) );
  HS65_LL_MUXI21X2 U16375 ( .D0(n15429), .D1(w3[12]), .S0(n15428), .Z(N469) );
  HS65_LL_MUXI21X2 U16376 ( .D0(w3[11]), .D1(n15431), .S0(n15430), .Z(N470) );
  HS65_LL_MUXI21X2 U16377 ( .D0(n15720), .D1(n15672), .S0(w3[10]), .Z(N471) );
  HS65_LL_MUXI21X2 U16378 ( .D0(n15433), .D1(w3[9]), .S0(n15432), .Z(N472) );
  HS65_LL_IVX2 U16379 ( .A(w3[8]), .Z(n15700) );
  HS65_LL_MUXI21X2 U16380 ( .D0(w3[8]), .D1(n15700), .S0(n15434), .Z(N473) );
  HS65_LL_MUXI21X2 U16381 ( .D0(n15436), .D1(n15435), .S0(w0[7]), .Z(N474) );
  HS65_LL_MUXI21X2 U16382 ( .D0(n15530), .D1(n15531), .S0(w0[6]), .Z(N475) );
  HS65_LL_IVX2 U16383 ( .A(n15521), .Z(n15437) );
  HS65_LL_MUXI21X2 U16384 ( .D0(n15437), .D1(n15521), .S0(w0[5]), .Z(N476) );
  HS65_LL_MUXI21X2 U16385 ( .D0(n15438), .D1(w0[4]), .S0(n15540), .Z(N477) );
  HS65_LL_MUXI21X2 U16386 ( .D0(w0[3]), .D1(n15440), .S0(n15439), .Z(N478) );
  HS65_LL_MUXI21X2 U16387 ( .D0(n15442), .D1(n15441), .S0(w0[1]), .Z(N480) );
  HS65_LL_MUXI21X2 U16388 ( .D0(n15550), .D1(n15551), .S0(w0[0]), .Z(N481) );
  HS65_LL_MUXI21X2 U16389 ( .D0(n15444), .D1(n15443), .S0(w1[7]), .Z(N482) );
  HS65_LL_IVX2 U16390 ( .A(n15445), .Z(n15446) );
  HS65_LL_MUXI21X2 U16391 ( .D0(n15446), .D1(n15445), .S0(w1[6]), .Z(N483) );
  HS65_LL_MUXI21X2 U16392 ( .D0(w1[4]), .D1(n15448), .S0(n15447), .Z(N485) );
  HS65_LL_MUXI21X2 U16393 ( .D0(w1[3]), .D1(n15450), .S0(n15449), .Z(N486) );
  HS65_LL_MUXI21X2 U16394 ( .D0(n15452), .D1(w1[1]), .S0(n15451), .Z(N488) );
  HS65_LL_MUXI21X2 U16395 ( .D0(n15454), .D1(n15453), .S0(w1[0]), .Z(N489) );
  HS65_LL_IVX2 U16396 ( .A(w2[7]), .Z(n15655) );
  HS65_LL_MUXI21X2 U16397 ( .D0(w2[7]), .D1(n15655), .S0(n15455), .Z(N490) );
  HS65_LL_IVX2 U16398 ( .A(w2[6]), .Z(n15646) );
  HS65_LL_MUXI21X2 U16399 ( .D0(n15646), .D1(w2[6]), .S0(n15587), .Z(N491) );
  HS65_LL_IVX2 U16400 ( .A(w2[5]), .Z(n15640) );
  HS65_LL_NAND4ABX3 U16401 ( .A(n15459), .B(n15458), .C(n15457), .D(n15456), 
        .Z(n15461) );
  HS65_LL_NAND4ABX3 U16402 ( .A(n15462), .B(n15461), .C(n15460), .D(n15474), 
        .Z(n15504) );
  HS65_LL_NAND4ABX3 U16403 ( .A(n15466), .B(n15465), .C(n15464), .D(n15463), 
        .Z(n15467) );
  HS65_LL_NOR4ABX2 U16404 ( .A(n15470), .B(n15469), .C(n15468), .D(n15467), 
        .Z(n15501) );
  HS65_LL_NOR4ABX2 U16405 ( .A(n15474), .B(n15473), .C(n15472), .D(n15471), 
        .Z(n15476) );
  HS65_LL_NAND4ABX3 U16406 ( .A(n15489), .B(n15477), .C(n15476), .D(n15475), 
        .Z(n15479) );
  HS65_LL_OAI13X1 U16407 ( .A(n15481), .B(n15480), .C(n15479), .D(n15478), .Z(
        n15499) );
  HS65_LL_NAND4ABX3 U16408 ( .A(n15485), .B(n15484), .C(n15483), .D(n15482), 
        .Z(n15488) );
  HS65_LL_NAND4ABX3 U16409 ( .A(n15489), .B(n15488), .C(n15487), .D(n15486), 
        .Z(n15492) );
  HS65_LL_NAND4ABX3 U16410 ( .A(n15493), .B(n15492), .C(n15491), .D(n15490), 
        .Z(n15495) );
  HS65_LL_OAI13X1 U16411 ( .A(n15497), .B(n15496), .C(n15495), .D(n15494), .Z(
        n15498) );
  HS65_LL_OAI112X1 U16412 ( .A(n15501), .B(n15500), .C(n15499), .D(n15498), 
        .Z(n15502) );
  HS65_LL_CBI4I6X2 U16413 ( .A(n15505), .B(n15504), .C(n15503), .D(n15502), 
        .Z(n15612) );
  HS65_LL_MUXI21X2 U16414 ( .D0(w2[5]), .D1(n15640), .S0(n15612), .Z(N492) );
  HS65_LL_MUXI21X2 U16415 ( .D0(n15507), .D1(w2[4]), .S0(n15506), .Z(N493) );
  HS65_LL_MUXI21X2 U16416 ( .D0(w2[3]), .D1(n15509), .S0(n15508), .Z(N494) );
  HS65_LL_IVX2 U16417 ( .A(w2[2]), .Z(n15634) );
  HS65_LL_MUXI21X2 U16418 ( .D0(w2[2]), .D1(n15634), .S0(n15510), .Z(N495) );
  HS65_LL_MUXI21X2 U16419 ( .D0(n15512), .D1(w2[1]), .S0(n15511), .Z(N496) );
  HS65_LL_IVX2 U16420 ( .A(w2[0]), .Z(n15628) );
  HS65_LL_IVX2 U16421 ( .A(n15561), .Z(n15562) );
  HS65_LL_MUXI21X2 U16422 ( .D0(w2[0]), .D1(n15628), .S0(n15562), .Z(N497) );
  HS65_LL_MUXI21X2 U16423 ( .D0(w3[7]), .D1(n15746), .S0(n15513), .Z(N498) );
  HS65_LL_MUXI21X2 U16424 ( .D0(w3[6]), .D1(n15737), .S0(n15682), .Z(N499) );
  HS65_LL_MUXI21X2 U16425 ( .D0(n15730), .D1(w3[5]), .S0(n15701), .Z(N500) );
  HS65_LL_MUXI21X2 U16426 ( .D0(w3[4]), .D1(n15515), .S0(n15514), .Z(N501) );
  HS65_LL_MUXI21X2 U16427 ( .D0(w3[3]), .D1(n15517), .S0(n15516), .Z(N502) );
  HS65_LL_MUXI21X2 U16428 ( .D0(w3[2]), .D1(n15723), .S0(n15518), .Z(N503) );
  HS65_LL_MUXI21X2 U16429 ( .D0(n15520), .D1(w3[1]), .S0(n15519), .Z(N504) );
  HS65_LL_MUXI21X2 U16430 ( .D0(w3[0]), .D1(n15717), .S0(n15657), .Z(N505) );
  HS65_LLS_XOR3X2 U16431 ( .A(w0[29]), .B(n15522), .C(n15521), .Z(n15525) );
  HS65_LLS_XOR3X2 U16432 ( .A(n15525), .B(n15524), .C(n15523), .Z(n15528) );
  HS65_LL_MUXI21X2 U16433 ( .D0(w0[29]), .D1(n15526), .S0(text_in_r[125]), .Z(
        n15527) );
  HS65_LL_MUXI21X2 U16434 ( .D0(n15528), .D1(n15527), .S0(n15688), .Z(N279) );
  HS65_LL_MUXI21X2 U16435 ( .D0(n15531), .D1(n15530), .S0(n15529), .Z(n15532)
         );
  HS65_LL_MUXI21X2 U16436 ( .D0(n15548), .D1(n15549), .S0(n15532), .Z(n15533)
         );
  HS65_LL_BDECNX4 U16437 ( .ZNP(w0[30]), .ZNN(n15534), .DNM1(n15533), .DN(
        text_in_r[126]), .NDBL(n15727), .Z(N280) );
  HS65_LLS_XOR3X2 U16438 ( .A(n15537), .B(n15536), .C(n15535), .Z(n15538) );
  HS65_LL_BDECNX4 U16439 ( .ZNP(w0[10]), .ZNN(n15539), .DNM1(n15538), .DN(
        text_in_r[106]), .NDBL(n15727), .Z(N244) );
  HS65_LL_MUXI21X2 U16440 ( .D0(n15541), .D1(w0[13]), .S0(text_in_r[109]), .Z(
        n15547) );
  HS65_LL_MUXI21X2 U16441 ( .D0(w0[13]), .D1(n15541), .S0(n15540), .Z(n15544)
         );
  HS65_LLS_XOR3X2 U16442 ( .A(n15544), .B(n15543), .C(n15542), .Z(n15546) );
  HS65_LL_MUX31X4 U16443 ( .D0(n15549), .D1(n15548), .D2(n15547), .S0(n15546), 
        .S1(n15545), .Z(N247) );
  HS65_LL_MUXI21X2 U16444 ( .D0(n15551), .D1(n15550), .S0(w0[1]), .Z(n15554)
         );
  HS65_LLS_XOR3X2 U16445 ( .A(n15554), .B(n15553), .C(n15552), .Z(n15555) );
  HS65_LLS_XOR3X2 U16446 ( .A(n15557), .B(n15556), .C(n15555), .Z(n15560) );
  HS65_LL_MUXI21X2 U16447 ( .D0(w0[1]), .D1(n15558), .S0(text_in_r[97]), .Z(
        n15559) );
  HS65_LL_MUXI21X2 U16448 ( .D0(n15560), .D1(n15559), .S0(n15688), .Z(N227) );
  HS65_LL_MUXI21X2 U16449 ( .D0(n15562), .D1(n15561), .S0(n15623), .Z(n15563)
         );
  HS65_LL_MUXI21X2 U16450 ( .D0(n15652), .D1(n15651), .S0(n15563), .Z(n15564)
         );
  HS65_LL_OAI21X2 U16451 ( .A(text_in_r[56]), .B(n11557), .C(n15564), .Z(
        n15565) );
  HS65_LL_MUXI21X2 U16452 ( .D0(w2[24]), .D1(n15566), .S0(n15565), .Z(N146) );
  HS65_LL_MUXI21X2 U16453 ( .D0(n15637), .D1(n15567), .S0(n15575), .Z(n15588)
         );
  HS65_LLS_XOR3X2 U16454 ( .A(n15612), .B(n15588), .C(w2[29]), .Z(n15570) );
  HS65_LLS_XOR3X2 U16455 ( .A(n15570), .B(n15569), .C(n15568), .Z(n15573) );
  HS65_LL_MUXI21X2 U16456 ( .D0(w2[29]), .D1(n15571), .S0(text_in_r[61]), .Z(
        n15572) );
  HS65_LL_MUXI21X2 U16457 ( .D0(n15573), .D1(n15572), .S0(n15734), .Z(N151) );
  HS65_LL_MUXI21X2 U16458 ( .D0(n15574), .D1(n15589), .S0(n15619), .Z(n15643)
         );
  HS65_LL_MUXI21X2 U16459 ( .D0(n15614), .D1(n15613), .S0(n15575), .Z(n15635)
         );
  HS65_LLS_XNOR3X2 U16460 ( .A(n15587), .B(n15643), .C(n15635), .Z(n15576) );
  HS65_LL_BDECNX4 U16461 ( .ZNP(w2[30]), .ZNN(n15577), .DNM1(n15576), .DN(
        text_in_r[62]), .NDBL(n15727), .Z(N152) );
  HS65_LLS_XOR3X2 U16462 ( .A(n15600), .B(n15579), .C(n15578), .Z(n15580) );
  HS65_LL_MUXI21X2 U16463 ( .D0(n15580), .D1(text_in_r[48]), .S0(n15734), .Z(
        n15581) );
  HS65_LL_MUXI21X2 U16464 ( .D0(w2[16]), .D1(n15582), .S0(n15581), .Z(N130) );
  HS65_LLS_XOR2X3 U16465 ( .A(n15612), .B(n15637), .Z(n15620) );
  HS65_LLS_XOR3X2 U16466 ( .A(n15583), .B(n15620), .C(n15614), .Z(n15584) );
  HS65_LL_MUXI21X2 U16467 ( .D0(n15584), .D1(text_in_r[53]), .S0(n15734), .Z(
        n15585) );
  HS65_LL_MUXI21X2 U16468 ( .D0(w2[21]), .D1(n15586), .S0(n15585), .Z(N135) );
  HS65_LLS_XOR2X3 U16469 ( .A(n15587), .B(n15641), .Z(n15647) );
  HS65_LLS_XOR3X2 U16470 ( .A(n15647), .B(n15589), .C(n15588), .Z(n15590) );
  HS65_LL_MUXI21X2 U16471 ( .D0(n15590), .D1(text_in_r[54]), .S0(n15734), .Z(
        n15591) );
  HS65_LL_MUXI21X2 U16472 ( .D0(w2[22]), .D1(n15592), .S0(n15591), .Z(N136) );
  HS65_LL_MUXI21X2 U16473 ( .D0(n15594), .D1(n15593), .S0(n15643), .Z(n15595)
         );
  HS65_LL_MUXI21X2 U16474 ( .D0(n15603), .D1(n15602), .S0(n15595), .Z(n15596)
         );
  HS65_LL_OAI21X2 U16475 ( .A(text_in_r[55]), .B(n11557), .C(n15596), .Z(
        n15597) );
  HS65_LL_MUXI21X2 U16476 ( .D0(w2[23]), .D1(n15598), .S0(n15597), .Z(N137) );
  HS65_LLS_XNOR2X3 U16477 ( .A(n15600), .B(n15599), .Z(n15601) );
  HS65_LL_MUXI21X2 U16478 ( .D0(n15603), .D1(n15602), .S0(n15601), .Z(n15604)
         );
  HS65_LL_OAI21X2 U16479 ( .A(text_in_r[40]), .B(n11557), .C(n15604), .Z(
        n15605) );
  HS65_LL_MUXI21X2 U16480 ( .D0(w2[8]), .D1(n15606), .S0(n15605), .Z(N114) );
  HS65_LL_IVX2 U16481 ( .A(w2[10]), .Z(n15611) );
  HS65_LLS_XOR3X2 U16482 ( .A(n15609), .B(n15608), .C(n15607), .Z(n15610) );
  HS65_LL_BDECNX4 U16483 ( .ZNP(w2[10]), .ZNN(n15611), .DNM1(n15610), .DN(
        text_in_r[42]), .NDBL(n15727), .Z(N116) );
  HS65_LL_MUXI21X2 U16484 ( .D0(n15614), .D1(n15613), .S0(n15612), .Z(n15642)
         );
  HS65_LLS_XOR3X2 U16485 ( .A(n15616), .B(n15642), .C(n15615), .Z(n15617) );
  HS65_LL_BDECNX4 U16486 ( .ZNP(w2[13]), .ZNN(n15618), .DNM1(n15617), .DN(
        text_in_r[45]), .NDBL(n15727), .Z(N119) );
  HS65_LLS_XOR3X2 U16487 ( .A(n15620), .B(n15647), .C(n15619), .Z(n15621) );
  HS65_LL_BDECNX4 U16488 ( .ZNP(w2[14]), .ZNN(n15622), .DNM1(n15621), .DN(
        text_in_r[46]), .NDBL(n15727), .Z(N120) );
  HS65_LLS_XOR3X2 U16489 ( .A(n15625), .B(n15624), .C(n15623), .Z(n15626) );
  HS65_LL_MUXI21X2 U16490 ( .D0(n15626), .D1(text_in_r[32]), .S0(n15734), .Z(
        n15627) );
  HS65_LL_MUXI21X2 U16491 ( .D0(w2[0]), .D1(n15628), .S0(n15627), .Z(N98) );
  HS65_LLS_XOR3X2 U16492 ( .A(n15631), .B(n15630), .C(n15629), .Z(n15632) );
  HS65_LL_MUXI21X2 U16493 ( .D0(n15632), .D1(text_in_r[34]), .S0(n15734), .Z(
        n15633) );
  HS65_LL_MUXI21X2 U16494 ( .D0(w2[2]), .D1(n15634), .S0(n15633), .Z(N100) );
  HS65_LLS_XOR3X2 U16495 ( .A(n15637), .B(n15636), .C(n15635), .Z(n15638) );
  HS65_LL_MUXI21X2 U16496 ( .D0(n15638), .D1(text_in_r[37]), .S0(n15734), .Z(
        n15639) );
  HS65_LL_MUXI21X2 U16497 ( .D0(w2[5]), .D1(n15640), .S0(n15639), .Z(N103) );
  HS65_LLS_XOR3X2 U16498 ( .A(n15643), .B(n15642), .C(n15641), .Z(n15644) );
  HS65_LL_MUXI21X2 U16499 ( .D0(n15644), .D1(text_in_r[38]), .S0(n15734), .Z(
        n15645) );
  HS65_LL_MUXI21X2 U16500 ( .D0(w2[6]), .D1(n15646), .S0(n15645), .Z(N104) );
  HS65_LL_MUXI21X2 U16501 ( .D0(n15649), .D1(n15648), .S0(n15647), .Z(n15650)
         );
  HS65_LL_MUXI21X2 U16502 ( .D0(n15652), .D1(n15651), .S0(n15650), .Z(n15653)
         );
  HS65_LL_OAI21X2 U16503 ( .A(text_in_r[39]), .B(n11557), .C(n15653), .Z(
        n15654) );
  HS65_LL_MUXI21X2 U16504 ( .D0(w2[7]), .D1(n15655), .S0(n15654), .Z(N105) );
  HS65_LL_MUXI21X2 U16505 ( .D0(n15657), .D1(n15656), .S0(n15712), .Z(n15658)
         );
  HS65_LL_MUXI21X2 U16506 ( .D0(n15743), .D1(n15742), .S0(n15658), .Z(n15659)
         );
  HS65_LL_OAI21X2 U16507 ( .A(text_in_r[24]), .B(n11557), .C(n15659), .Z(
        n15660) );
  HS65_LL_MUXI21X2 U16508 ( .D0(w3[24]), .D1(n15661), .S0(n15660), .Z(N82) );
  HS65_LL_MUXI21X2 U16509 ( .D0(n15683), .D1(n15663), .S0(n15662), .Z(n15732)
         );
  HS65_LL_MUXI21X2 U16510 ( .D0(n15703), .D1(n15702), .S0(n15664), .Z(n15724)
         );
  HS65_LLS_XOR3X2 U16511 ( .A(n15682), .B(n15732), .C(n15724), .Z(n15665) );
  HS65_LL_BDECNX4 U16512 ( .ZNP(w3[30]), .ZNN(n15666), .DNM1(n15665), .DN(
        text_in_r[30]), .NDBL(n15727), .Z(N88) );
  HS65_LLS_XOR3X2 U16513 ( .A(n15692), .B(n15668), .C(n15667), .Z(n15669) );
  HS65_LL_MUXI21X2 U16514 ( .D0(n15669), .D1(text_in_r[16]), .S0(n15734), .Z(
        n15670) );
  HS65_LL_MUXI21X2 U16515 ( .D0(w3[16]), .D1(n15671), .S0(n15670), .Z(N66) );
  HS65_LLS_XOR3X2 U16516 ( .A(n15674), .B(n15673), .C(n15672), .Z(n15675) );
  HS65_LL_MUXI21X2 U16517 ( .D0(n15675), .D1(text_in_r[18]), .S0(n15734), .Z(
        n15676) );
  HS65_LL_MUXI21X2 U16518 ( .D0(w3[18]), .D1(n15785), .S0(n15676), .Z(N68) );
  HS65_LLS_XOR2X3 U16519 ( .A(n15701), .B(n15677), .Z(n15709) );
  HS65_LLS_XOR3X2 U16520 ( .A(n15678), .B(n15709), .C(n15703), .Z(n15679) );
  HS65_LL_MUXI21X2 U16521 ( .D0(n15679), .D1(text_in_r[21]), .S0(n15727), .Z(
        n15680) );
  HS65_LL_MUXI21X2 U16522 ( .D0(w3[21]), .D1(n15681), .S0(n15680), .Z(N71) );
  HS65_LLS_XOR2X3 U16523 ( .A(n15733), .B(n15682), .Z(n15738) );
  HS65_LLS_XOR3X2 U16524 ( .A(n15738), .B(n15684), .C(n15683), .Z(n15685) );
  HS65_LL_MUXI21X2 U16525 ( .D0(n15685), .D1(text_in_r[22]), .S0(n15734), .Z(
        n15686) );
  HS65_LL_MUXI21X2 U16526 ( .D0(w3[22]), .D1(n15687), .S0(n15686), .Z(N72) );
  HS65_LLS_XOR3X2 U16527 ( .A(n15739), .B(n15732), .C(n15713), .Z(n15689) );
  HS65_LL_MUXI21X2 U16528 ( .D0(n15689), .D1(text_in_r[23]), .S0(n15688), .Z(
        n15690) );
  HS65_LL_MUXI21X2 U16529 ( .D0(w3[23]), .D1(n15691), .S0(n15690), .Z(N73) );
  HS65_LL_MUX21I1X3 U16530 ( .D0(n15693), .D1(n15693), .S0(n15692), .Z(n15694)
         );
  HS65_LL_MUX21X4 U16531 ( .D0(n15696), .D1(n15695), .S0(n15694), .Z(n15697)
         );
  HS65_LL_AOI12X2 U16532 ( .A(n15698), .B(text_in_r[8]), .C(n15697), .Z(n15699) );
  HS65_LL_MUXI21X2 U16533 ( .D0(w3[8]), .D1(n15700), .S0(n15699), .Z(N50) );
  HS65_LL_MUXI21X2 U16534 ( .D0(n15703), .D1(n15702), .S0(n15701), .Z(n15731)
         );
  HS65_LLS_XOR3X2 U16535 ( .A(n15705), .B(n15704), .C(n15731), .Z(n15706) );
  HS65_LL_BDECNX4 U16536 ( .ZNP(w3[13]), .ZNN(n15707), .DNM1(n15706), .DN(
        text_in_r[13]), .NDBL(n15727), .Z(N55) );
  HS65_LLS_XOR3X2 U16537 ( .A(n15709), .B(n15738), .C(n15708), .Z(n15710) );
  HS65_LL_BDECNX4 U16538 ( .ZNP(w3[14]), .ZNN(n15711), .DNM1(n15710), .DN(
        text_in_r[14]), .NDBL(n15727), .Z(N56) );
  HS65_LLS_XOR3X2 U16539 ( .A(n15714), .B(n15713), .C(n15712), .Z(n15715) );
  HS65_LL_MUXI21X2 U16540 ( .D0(n15715), .D1(text_in_r[0]), .S0(n15727), .Z(
        n15716) );
  HS65_LL_MUXI21X2 U16541 ( .D0(w3[0]), .D1(n15717), .S0(n15716), .Z(N34) );
  HS65_LLS_XOR3X2 U16542 ( .A(n15720), .B(n15719), .C(n15718), .Z(n15721) );
  HS65_LL_MUXI21X2 U16543 ( .D0(n15721), .D1(text_in_r[2]), .S0(n15727), .Z(
        n15722) );
  HS65_LL_MUXI21X2 U16544 ( .D0(w3[2]), .D1(n15723), .S0(n15722), .Z(N36) );
  HS65_LLS_XOR3X2 U16545 ( .A(n15726), .B(n15725), .C(n15724), .Z(n15728) );
  HS65_LL_MUXI21X2 U16546 ( .D0(n15728), .D1(text_in_r[5]), .S0(n15727), .Z(
        n15729) );
  HS65_LL_MUXI21X2 U16547 ( .D0(w3[5]), .D1(n15730), .S0(n15729), .Z(N39) );
  HS65_LLS_XOR3X2 U16548 ( .A(n15733), .B(n15732), .C(n15731), .Z(n15735) );
  HS65_LL_MUXI21X2 U16549 ( .D0(n15735), .D1(text_in_r[6]), .S0(n15734), .Z(
        n15736) );
  HS65_LL_MUXI21X2 U16550 ( .D0(w3[6]), .D1(n15737), .S0(n15736), .Z(N40) );
  HS65_LL_MUXI21X2 U16551 ( .D0(n15740), .D1(n15739), .S0(n15738), .Z(n15741)
         );
  HS65_LL_MUXI21X2 U16552 ( .D0(n15743), .D1(n15742), .S0(n15741), .Z(n15744)
         );
  HS65_LL_OAI21X2 U16553 ( .A(text_in_r[7]), .B(n11557), .C(n15744), .Z(n15745) );
  HS65_LL_MUXI21X2 U16554 ( .D0(w3[7]), .D1(n15746), .S0(n15745), .Z(N41) );
  HS65_LL_NOR2AX3 U16555 ( .A(n15748), .B(n15747), .Z(\u0/r0/N76 ) );
  HS65_LL_MUXI21X2 U16556 ( .D0(key[0]), .D1(w3[0]), .S0(n15844), .Z(n15750)
         );
  HS65_LL_MUXI21X2 U16557 ( .D0(n15750), .D1(w3[0]), .S0(n15749), .Z(\u0/N240 ) );
  HS65_LL_MUXI21X2 U16558 ( .D0(key[1]), .D1(w3[1]), .S0(n15844), .Z(n15752)
         );
  HS65_LL_MUXI21X2 U16559 ( .D0(n15752), .D1(w3[1]), .S0(n15751), .Z(\u0/N241 ) );
  HS65_LL_MUXI21X2 U16560 ( .D0(key[2]), .D1(w3[2]), .S0(n15844), .Z(n15754)
         );
  HS65_LL_MUXI21X2 U16561 ( .D0(n15754), .D1(w3[2]), .S0(n15753), .Z(\u0/N242 ) );
  HS65_LL_MUXI21X2 U16562 ( .D0(key[3]), .D1(w3[3]), .S0(n15844), .Z(n15756)
         );
  HS65_LL_MUXI21X2 U16563 ( .D0(n15756), .D1(w3[3]), .S0(n15755), .Z(\u0/N243 ) );
  HS65_LL_MUXI21X2 U16564 ( .D0(key[4]), .D1(w3[4]), .S0(n15806), .Z(n15758)
         );
  HS65_LL_MUXI21X2 U16565 ( .D0(n15758), .D1(w3[4]), .S0(n15757), .Z(\u0/N244 ) );
  HS65_LL_MUXI21X2 U16566 ( .D0(key[5]), .D1(w3[5]), .S0(n15806), .Z(n15760)
         );
  HS65_LL_MUXI21X2 U16567 ( .D0(n15760), .D1(w3[5]), .S0(n15759), .Z(\u0/N245 ) );
  HS65_LL_MUXI21X2 U16568 ( .D0(key[6]), .D1(w3[6]), .S0(n15806), .Z(n15762)
         );
  HS65_LL_MUXI21X2 U16569 ( .D0(n15762), .D1(w3[6]), .S0(n15761), .Z(\u0/N246 ) );
  HS65_LL_MUXI21X2 U16570 ( .D0(key[7]), .D1(w3[7]), .S0(n15843), .Z(n15764)
         );
  HS65_LL_MUXI21X2 U16571 ( .D0(n15764), .D1(w3[7]), .S0(n15763), .Z(\u0/N247 ) );
  HS65_LL_MUXI21X2 U16572 ( .D0(key[8]), .D1(w3[8]), .S0(n15843), .Z(n15766)
         );
  HS65_LL_MUXI21X2 U16573 ( .D0(n15766), .D1(w3[8]), .S0(n15765), .Z(\u0/N248 ) );
  HS65_LL_MUXI21X2 U16574 ( .D0(key[9]), .D1(w3[9]), .S0(n15843), .Z(n15768)
         );
  HS65_LL_MUXI21X2 U16575 ( .D0(n15768), .D1(w3[9]), .S0(n15767), .Z(\u0/N249 ) );
  HS65_LL_MUXI21X2 U16576 ( .D0(key[10]), .D1(w3[10]), .S0(n15843), .Z(n15770)
         );
  HS65_LL_MUXI21X2 U16577 ( .D0(n15770), .D1(w3[10]), .S0(n15769), .Z(
        \u0/N250 ) );
  HS65_LL_MUXI21X2 U16578 ( .D0(key[11]), .D1(w3[11]), .S0(n15843), .Z(n15772)
         );
  HS65_LL_MUXI21X2 U16579 ( .D0(n15772), .D1(w3[11]), .S0(n15771), .Z(
        \u0/N251 ) );
  HS65_LL_MUXI21X2 U16580 ( .D0(key[12]), .D1(w3[12]), .S0(n15843), .Z(n15774)
         );
  HS65_LL_MUXI21X2 U16581 ( .D0(n15774), .D1(w3[12]), .S0(n15773), .Z(
        \u0/N252 ) );
  HS65_LL_MUXI21X2 U16582 ( .D0(key[14]), .D1(w3[14]), .S0(n15843), .Z(n15776)
         );
  HS65_LL_MUXI21X2 U16583 ( .D0(n15776), .D1(w3[14]), .S0(n15775), .Z(
        \u0/N254 ) );
  HS65_LL_MUXI21X2 U16584 ( .D0(key[15]), .D1(w3[15]), .S0(n15843), .Z(n15778)
         );
  HS65_LL_MUXI21X2 U16585 ( .D0(n15778), .D1(w3[15]), .S0(n15777), .Z(
        \u0/N255 ) );
  HS65_LL_MUXI21X2 U16586 ( .D0(key[16]), .D1(w3[16]), .S0(n15843), .Z(n15780)
         );
  HS65_LL_MUXI21X2 U16587 ( .D0(n15780), .D1(w3[16]), .S0(n15779), .Z(
        \u0/N256 ) );
  HS65_LL_MUXI21X2 U16588 ( .D0(key[17]), .D1(w3[17]), .S0(n15844), .Z(n15782)
         );
  HS65_LL_MUXI21X2 U16589 ( .D0(n15782), .D1(w3[17]), .S0(n15781), .Z(
        \u0/N257 ) );
  HS65_LL_MUX31X4 U16590 ( .D0(n15785), .D1(w3[18]), .D2(key[18]), .S0(n15784), 
        .S1(n15783), .Z(\u0/N258 ) );
  HS65_LL_MUXI21X2 U16591 ( .D0(key[19]), .D1(w3[19]), .S0(n15844), .Z(n15787)
         );
  HS65_LL_MUXI21X2 U16592 ( .D0(n15787), .D1(w3[19]), .S0(n15786), .Z(
        \u0/N259 ) );
  HS65_LL_MUXI21X2 U16593 ( .D0(key[20]), .D1(w3[20]), .S0(n15844), .Z(n15789)
         );
  HS65_LL_MUXI21X2 U16594 ( .D0(n15789), .D1(w3[20]), .S0(n15788), .Z(
        \u0/N260 ) );
  HS65_LL_MUXI21X2 U16595 ( .D0(key[21]), .D1(w3[21]), .S0(n15844), .Z(n15791)
         );
  HS65_LL_MUXI21X2 U16596 ( .D0(n15791), .D1(w3[21]), .S0(n15790), .Z(
        \u0/N261 ) );
  HS65_LL_MUXI21X2 U16597 ( .D0(key[22]), .D1(w3[22]), .S0(n15844), .Z(n15793)
         );
  HS65_LL_MUXI21X2 U16598 ( .D0(n15793), .D1(w3[22]), .S0(n15792), .Z(
        \u0/N262 ) );
  HS65_LL_MUXI21X2 U16599 ( .D0(key[23]), .D1(w3[23]), .S0(n15806), .Z(n15795)
         );
  HS65_LL_MUXI21X2 U16600 ( .D0(n15795), .D1(w3[23]), .S0(n15794), .Z(
        \u0/N263 ) );
  HS65_LL_MUXI21X2 U16601 ( .D0(key[24]), .D1(w3[24]), .S0(n15844), .Z(n15797)
         );
  HS65_LL_MUXI21X2 U16602 ( .D0(n15797), .D1(w3[24]), .S0(n15796), .Z(
        \u0/N264 ) );
  HS65_LL_MUXI21X2 U16603 ( .D0(key[26]), .D1(w3[26]), .S0(n15806), .Z(n15799)
         );
  HS65_LL_MUXI21X2 U16604 ( .D0(n15799), .D1(w3[26]), .S0(n15798), .Z(
        \u0/N266 ) );
  HS65_LL_MUXI21X2 U16605 ( .D0(key[27]), .D1(w3[27]), .S0(n15806), .Z(n15801)
         );
  HS65_LL_MUXI21X2 U16606 ( .D0(n15801), .D1(w3[27]), .S0(n15800), .Z(
        \u0/N267 ) );
  HS65_LL_MUXI21X2 U16607 ( .D0(key[28]), .D1(w3[28]), .S0(n15844), .Z(n15803)
         );
  HS65_LL_MUXI21X2 U16608 ( .D0(n15803), .D1(w3[28]), .S0(n15802), .Z(
        \u0/N268 ) );
  HS65_LL_MUXI21X2 U16609 ( .D0(key[30]), .D1(w3[30]), .S0(n15806), .Z(n15805)
         );
  HS65_LL_MUXI21X2 U16610 ( .D0(n15805), .D1(w3[30]), .S0(n15804), .Z(
        \u0/N270 ) );
  HS65_LL_MUXI21X2 U16611 ( .D0(key[31]), .D1(w3[31]), .S0(n15806), .Z(n15808)
         );
  HS65_LL_MUXI21X2 U16612 ( .D0(n15808), .D1(w3[31]), .S0(n15807), .Z(
        \u0/N271 ) );
  HS65_LL_MUX21X4 U16613 ( .D0(n15809), .D1(key[64]), .S0(n15826), .Z(
        \u0/N108 ) );
  HS65_LL_MUX21X4 U16614 ( .D0(n15810), .D1(key[65]), .S0(n15826), .Z(
        \u0/N109 ) );
  HS65_LL_MUX21X4 U16615 ( .D0(n15811), .D1(key[66]), .S0(n15826), .Z(
        \u0/N110 ) );
  HS65_LL_MUX21X4 U16616 ( .D0(n15812), .D1(key[67]), .S0(n15826), .Z(
        \u0/N111 ) );
  HS65_LL_MUX21X4 U16617 ( .D0(n15813), .D1(key[68]), .S0(n15826), .Z(
        \u0/N112 ) );
  HS65_LL_MUX21X4 U16618 ( .D0(n15814), .D1(key[69]), .S0(n15826), .Z(
        \u0/N113 ) );
  HS65_LL_MUX21X4 U16619 ( .D0(n15815), .D1(key[70]), .S0(n15826), .Z(
        \u0/N114 ) );
  HS65_LL_MUX21X4 U16620 ( .D0(n15816), .D1(key[71]), .S0(n15826), .Z(
        \u0/N115 ) );
  HS65_LL_IVX4 U16621 ( .A(n15844), .Z(n15839) );
  HS65_LL_MUX21X4 U16622 ( .D0(n15817), .D1(key[72]), .S0(n15839), .Z(
        \u0/N116 ) );
  HS65_LL_MUX21X4 U16623 ( .D0(n15818), .D1(key[73]), .S0(n15826), .Z(
        \u0/N117 ) );
  HS65_LL_MUX21X4 U16624 ( .D0(n15819), .D1(key[74]), .S0(n15826), .Z(
        \u0/N118 ) );
  HS65_LL_MUX21X4 U16625 ( .D0(n15820), .D1(key[75]), .S0(n15826), .Z(
        \u0/N119 ) );
  HS65_LL_MUX21X4 U16626 ( .D0(n15821), .D1(key[76]), .S0(n15826), .Z(
        \u0/N120 ) );
  HS65_LL_MUX21X4 U16627 ( .D0(n15822), .D1(key[78]), .S0(n15839), .Z(
        \u0/N122 ) );
  HS65_LL_MUX21X4 U16628 ( .D0(n15823), .D1(key[79]), .S0(n15826), .Z(
        \u0/N123 ) );
  HS65_LL_MUX21X4 U16629 ( .D0(n15824), .D1(key[80]), .S0(n15826), .Z(
        \u0/N124 ) );
  HS65_LL_MUX21X4 U16630 ( .D0(n15825), .D1(key[81]), .S0(n15839), .Z(
        \u0/N125 ) );
  HS65_LL_MUX21X4 U16631 ( .D0(n15827), .D1(key[82]), .S0(n15826), .Z(
        \u0/N126 ) );
  HS65_LL_MUX21X4 U16632 ( .D0(n15828), .D1(key[83]), .S0(n15839), .Z(
        \u0/N127 ) );
  HS65_LL_MUX21X4 U16633 ( .D0(n15829), .D1(key[84]), .S0(n15839), .Z(
        \u0/N128 ) );
  HS65_LL_MUX21X4 U16634 ( .D0(n15830), .D1(key[85]), .S0(n15839), .Z(
        \u0/N129 ) );
  HS65_LL_MUX21X4 U16635 ( .D0(n15831), .D1(key[86]), .S0(n15839), .Z(
        \u0/N130 ) );
  HS65_LL_MUX21X4 U16636 ( .D0(n15832), .D1(key[87]), .S0(n15839), .Z(
        \u0/N131 ) );
  HS65_LL_MUX21X4 U16637 ( .D0(n15833), .D1(key[88]), .S0(n15839), .Z(
        \u0/N132 ) );
  HS65_LL_MUX21X4 U16638 ( .D0(n15834), .D1(key[90]), .S0(n15839), .Z(
        \u0/N134 ) );
  HS65_LL_MUX21X4 U16639 ( .D0(n15835), .D1(key[91]), .S0(n15839), .Z(
        \u0/N135 ) );
  HS65_LL_MUX21X4 U16640 ( .D0(n15836), .D1(key[92]), .S0(n15839), .Z(
        \u0/N136 ) );
  HS65_LL_MUX21X4 U16641 ( .D0(n15837), .D1(key[94]), .S0(n15839), .Z(
        \u0/N138 ) );
  HS65_LL_MUX21X4 U16642 ( .D0(n15838), .D1(key[95]), .S0(n15839), .Z(
        \u0/N139 ) );
  HS65_LL_MUX21X4 U16643 ( .D0(n15840), .D1(key[127]), .S0(n15839), .Z(
        \u0/N73 ) );
  HS65_LL_AND2X4 U16644 ( .A(n15841), .B(n7668), .Z(n1) );
endmodule

