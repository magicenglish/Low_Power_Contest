
module c5315 ( N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, 
        N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, 
        N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
        N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
        N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, 
        N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, 
        N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, 
        N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
        N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, 
        N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, 
        N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, 
        N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, 
        N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
        N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, 
        N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, 
        N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, 
        N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, 
        N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, 
        N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, 
        N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, 
        N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, 
        N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, 
        N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, 
        N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, 
        N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, 
        N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, 
        N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128 );
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37,
         N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79,
         N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106,
         N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136,
         N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164,
         N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197,
         N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234,
         N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273,
         N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
         N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358,
         N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422,
         N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545,
         N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583,
         N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610,
         N613, N616, N619, N625, N631;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060,
         N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
         N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737,
         N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716,
         N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449,
         N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476,
         N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520,
         N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
         N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754,
         N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
         N8124, N8127, N8128;
  wire   N0, n1008, N6648, N6927, N4275, n1009, N1137, N1141, n485, n486, n488,
         n490, n492, n494, n496, n498, n500, n502, n504, n506, n508, n510,
         n512, N6926, n514, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n757, n758,
         n759, n760, n761, n762, n763, n764, n767, n768, n769, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n789, n791, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, N6643, N2527, N709, N2309;
  assign N1972 = N0;
  assign N6641 = N6648;
  assign N6925 = N6927;
  assign N4278 = N4275;
  assign N1143 = N1137;
  assign N1142 = N1137;
  assign N2584 = N1141;
  assign N6924 = N6926;
  assign N6646 = N6643;
  assign N3604 = N2527;
  assign N2142 = N709;
  assign N3360 = N2309;
  assign N3359 = N2309;
  assign N3358 = N2309;
  assign N3357 = N2309;

  HS65_LL_MX41X14 U544 ( .D0(n718), .S0(n973), .D1(n719), .S1(n974), .D2(n971), 
        .S2(N20), .D3(n972), .S3(N76), .Z(N7516) );
  HS65_LL_MX41X14 U545 ( .D0(n718), .S0(n968), .D1(n719), .S1(n967), .D2(n966), 
        .S2(N20), .D3(n965), .S3(N76), .Z(N7520) );
  HS65_LL_AO222X9 U546 ( .A(n918), .B(n516), .C(n806), .D(N114), .E(n921), .F(
        n885), .Z(n522) );
  HS65_LL_AOI21X2 U547 ( .A(n746), .B(n745), .C(n744), .Z(n747) );
  HS65_LL_NAND3X5 U548 ( .A(n675), .B(n674), .C(n673), .Z(n901) );
  HS65_LL_OAI222X2 U549 ( .A(n823), .B(n731), .C(n734), .D(n655), .E(n882), 
        .F(n654), .Z(n669) );
  HS65_LL_IVX35 U550 ( .A(n486), .Z(N7465) );
  HS65_LL_MUXI21X5 U551 ( .D0(n553), .D1(n552), .S0(N566), .Z(n554) );
  HS65_LLS_XNOR2X6 U552 ( .A(n566), .B(n540), .Z(n553) );
  HS65_LL_PAOI2X1 U553 ( .A(n861), .B(n566), .P(n696), .Z(n948) );
  HS65_LL_OAI12X3 U554 ( .A(n833), .B(N514), .C(n684), .Z(n713) );
  HS65_LL_AOI12X12 U555 ( .A(n562), .B(n739), .C(n559), .Z(n794) );
  HS65_LL_IVX2 U556 ( .A(n908), .Z(n485) );
  HS65_LL_NAND2X7 U557 ( .A(n805), .B(n804), .Z(n907) );
  HS65_LL_IVX18 U558 ( .A(n969), .Z(N7699) );
  HS65_LL_IVX9 U559 ( .A(n1009), .Z(n486) );
  HS65_LL_AOI12X3 U560 ( .A(n806), .B(N52), .C(n689), .Z(n1009) );
  HS65_LL_IVX2 U561 ( .A(n1008), .Z(n488) );
  HS65_LL_IVX18 U562 ( .A(n488), .Z(N2054) );
  HS65_LL_NOR2AX3 U563 ( .A(N136), .B(N1066), .Z(n1008) );
  HS65_LL_AND2X18 U564 ( .A(n521), .B(n527), .Z(N5388) );
  HS65_LL_IVX2 U565 ( .A(n668), .Z(n490) );
  HS65_LL_IVX18 U566 ( .A(n490), .Z(N7449) );
  HS65_LL_IVX2 U567 ( .A(n751), .Z(n492) );
  HS65_LL_IVX18 U568 ( .A(n492), .Z(N7607) );
  HS65_LL_IVX2 U569 ( .A(n754), .Z(n494) );
  HS65_LL_IVX18 U570 ( .A(n494), .Z(N7606) );
  HS65_LL_IVX2 U571 ( .A(n755), .Z(n496) );
  HS65_LL_IVX18 U572 ( .A(n496), .Z(N7605) );
  HS65_LL_IVX2 U573 ( .A(n662), .Z(n498) );
  HS65_LL_IVX18 U574 ( .A(n498), .Z(N7511) );
  HS65_LL_IVX2 U575 ( .A(n757), .Z(n500) );
  HS65_LL_IVX18 U576 ( .A(n500), .Z(N7601) );
  HS65_LL_IVX2 U577 ( .A(n666), .Z(n502) );
  HS65_LL_IVX18 U578 ( .A(n502), .Z(N7506) );
  HS65_LL_IVX2 U579 ( .A(n735), .Z(n504) );
  HS65_LL_IVX18 U580 ( .A(n504), .Z(N7522) );
  HS65_LL_IVX2 U581 ( .A(n711), .Z(n506) );
  HS65_LL_IVX18 U582 ( .A(n506), .Z(N7521) );
  HS65_LL_MX41X14 U583 ( .D0(n669), .S0(n968), .D1(n832), .S1(n967), .D2(n966), 
        .S2(N61), .D3(n965), .S3(N11), .Z(N7469) );
  HS65_LL_IVX2 U584 ( .A(n819), .Z(n508) );
  HS65_LL_IVX18 U585 ( .A(n508), .Z(N5240) );
  HS65_LL_NOR4ABX2 U586 ( .A(n818), .B(n817), .C(n816), .D(n815), .Z(n819) );
  HS65_LL_IVX2 U587 ( .A(n526), .Z(n510) );
  HS65_LL_IVX18 U588 ( .A(n510), .Z(N4272) );
  HS65_LL_OAI212X3 U589 ( .A(N588), .B(N86), .C(n947), .D(N87), .E(n906), .Z(
        n526) );
  HS65_LL_IVX2 U590 ( .A(n955), .Z(n512) );
  HS65_LL_IVX27 U591 ( .A(n512), .Z(N6926) );
  HS65_LL_OAI21X3 U592 ( .A(n954), .B(n953), .C(n952), .Z(n955) );
  HS65_LL_AOI12X2 U593 ( .A(N566), .B(n937), .C(n948), .Z(n567) );
  HS65_LL_AOI12X2 U594 ( .A(n748), .B(n672), .C(n943), .Z(n627) );
  HS65_LL_NAND2X2 U595 ( .A(n885), .B(n880), .Z(n639) );
  HS65_LL_MUXI21X2 U596 ( .D0(N233), .D1(N226), .S0(n853), .Z(n865) );
  HS65_LL_BFX9 U597 ( .A(n727), .Z(n514) );
  HS65_LL_MUXI41X2 U598 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n953), .S1(N206), .Z(n679) );
  HS65_LL_OAI21X2 U599 ( .A(n743), .B(n742), .C(n741), .Z(n928) );
  HS65_LL_OAI21X2 U600 ( .A(N400), .B(n705), .C(n704), .Z(n930) );
  HS65_LL_AOI12X2 U601 ( .A(N54), .B(n835), .C(n723), .Z(n823) );
  HS65_LL_IVX18 U602 ( .A(n528), .Z(N7701) );
  HS65_LL_AOI12X6 U603 ( .A(n937), .B(N4), .C(n948), .Z(n795) );
  HS65_LL_MUXI21X5 U604 ( .D0(n642), .D1(n960), .S0(n663), .Z(n644) );
  HS65_LL_AO12X18 U605 ( .A(n671), .B(N54), .C(n942), .Z(n745) );
  HS65_LLS_XNOR2X6 U606 ( .A(n677), .B(n558), .Z(n569) );
  HS65_LL_AOI12X6 U607 ( .A(n533), .B(n706), .C(n691), .Z(n566) );
  HS65_LL_MUXI21X10 U608 ( .D0(N358), .D1(N351), .S0(n842), .Z(n839) );
  HS65_LL_XOR3X9 U609 ( .A(n551), .B(n550), .C(n549), .Z(n552) );
  HS65_LL_MUXI21X5 U610 ( .D0(n740), .D1(n739), .S0(n738), .Z(n916) );
  HS65_LL_BFX27 U611 ( .A(n645), .Z(N8127) );
  HS65_LL_IVX9 U612 ( .A(N7465), .Z(n767) );
  HS65_LL_MX41X7 U613 ( .D0(n719), .S0(n959), .D1(n718), .S1(n958), .D2(n957), 
        .S2(N146), .D3(n956), .S3(N149), .Z(n751) );
  HS65_LL_IVX2 U614 ( .A(n907), .Z(n908) );
  HS65_LL_OAI12X3 U615 ( .A(n805), .B(n804), .C(n907), .Z(n826) );
  HS65_LL_NAND2X4 U616 ( .A(n516), .B(n915), .Z(n760) );
  HS65_LL_NAND2X4 U617 ( .A(n516), .B(n824), .Z(n673) );
  HS65_LL_MX41X7 U618 ( .D0(n769), .S0(n968), .D1(n768), .S1(n967), .D2(n966), 
        .S2(N70), .D3(n965), .S3(N67), .Z(n735) );
  HS65_LL_AOI22X3 U619 ( .A(n951), .B(n950), .C(n949), .D(n948), .Z(n952) );
  HS65_LL_IVX4 U620 ( .A(N7473), .Z(n768) );
  HS65_LL_AOI21X2 U621 ( .A(n671), .B(N583), .C(n942), .Z(n623) );
  HS65_LL_IVX4 U622 ( .A(N7363), .Z(n769) );
  HS65_LL_NOR3X3 U623 ( .A(n936), .B(n935), .C(n934), .Z(n949) );
  HS65_LL_OAI12X3 U624 ( .A(n653), .B(n739), .C(n935), .Z(n556) );
  HS65_LL_NOR3X1 U625 ( .A(N6877), .B(N1155), .C(N1152), .Z(n875) );
  HS65_LL_NAND2X4 U626 ( .A(n653), .B(n739), .Z(n935) );
  HS65_LL_NOR2X3 U627 ( .A(n723), .B(n822), .Z(n722) );
  HS65_LL_NOR2X3 U628 ( .A(n562), .B(n737), .Z(n653) );
  HS65_LL_NAND2X4 U629 ( .A(n615), .B(n746), .Z(n672) );
  HS65_LL_NAND2X4 U630 ( .A(N490), .B(n611), .Z(n615) );
  HS65_LL_IVX4 U631 ( .A(n869), .Z(n868) );
  HS65_LL_IVX4 U632 ( .A(n806), .Z(n734) );
  HS65_LL_IVX9 U633 ( .A(N2139), .Z(n665) );
  HS65_LL_NAND2X7 U634 ( .A(n888), .B(n886), .Z(n882) );
  HS65_LL_NAND2X5 U635 ( .A(n888), .B(N619), .Z(n731) );
  HS65_LL_IVX9 U636 ( .A(N625), .Z(n888) );
  HS65_LL_IVX4 U637 ( .A(N446), .Z(n953) );
  HS65_LL_IVX4 U638 ( .A(N435), .Z(n696) );
  HS65_LL_IVX4 U639 ( .A(N503), .Z(n688) );
  HS65_LL_IVX4 U640 ( .A(N571), .Z(n663) );
  HS65_LL_IVX9 U641 ( .A(n975), .Z(n642) );
  HS65_LL_AOI12X4 U642 ( .A(n516), .B(n887), .C(n574), .Z(n585) );
  HS65_LL_AOI22X1 U643 ( .A(N120), .B(N625), .C(N619), .D(n878), .Z(n879) );
  HS65_LL_AO222X9 U644 ( .A(n826), .B(n516), .C(n806), .D(N121), .E(n885), .F(
        n811), .Z(n807) );
  HS65_LL_AOI21X4 U645 ( .A(n516), .B(n877), .C(n641), .Z(n960) );
  HS65_LL_NAND2X5 U646 ( .A(n717), .B(n529), .Z(n718) );
  HS65_LL_NAND2X4 U647 ( .A(n547), .B(n546), .Z(n550) );
  HS65_LL_MX41X7 U648 ( .D0(n768), .S0(n964), .D1(n769), .S1(n963), .D2(n962), 
        .S2(N158), .D3(n961), .S3(N188), .Z(n757) );
  HS65_LL_MX41X7 U649 ( .D0(n523), .S0(n959), .D1(n524), .S1(n958), .D2(n957), 
        .S2(N152), .D3(n956), .S3(N155), .Z(n754) );
  HS65_LL_MX41X7 U650 ( .D0(n524), .S0(n968), .D1(n523), .S1(n967), .D2(n966), 
        .S2(N17), .D3(n965), .S3(N73), .Z(n711) );
  HS65_LL_MX41X7 U651 ( .D0(n768), .S0(n959), .D1(n769), .S1(n958), .D2(n957), 
        .S2(N158), .D3(n956), .S3(N188), .Z(n755) );
  HS65_LLS_XNOR2X3 U652 ( .A(n607), .B(n606), .Z(n609) );
  HS65_LL_NOR2X6 U653 ( .A(n695), .B(n565), .Z(n937) );
  HS65_LLS_XNOR2X3 U654 ( .A(n597), .B(n596), .Z(n607) );
  HS65_LL_NAND2X4 U655 ( .A(n640), .B(n639), .Z(n641) );
  HS65_LL_NOR2X3 U656 ( .A(n702), .B(n701), .Z(n681) );
  HS65_LL_MX41X7 U657 ( .D0(n832), .S0(n959), .D1(n669), .S1(n958), .D2(n957), 
        .S2(N185), .D3(n956), .S3(N182), .Z(n662) );
  HS65_LL_NOR2X6 U658 ( .A(n730), .B(n660), .Z(n707) );
  HS65_LL_MX41X7 U659 ( .D0(n669), .S0(n973), .D1(n832), .S1(n974), .D2(n971), 
        .S2(N61), .D3(n972), .S3(N11), .Z(n668) );
  HS65_LL_NAND2X7 U660 ( .A(n534), .B(n536), .Z(n706) );
  HS65_LL_MX41X7 U661 ( .D0(n832), .S0(n964), .D1(n669), .S1(n963), .D2(n962), 
        .S2(N185), .D3(n961), .S3(N182), .Z(n666) );
  HS65_LL_OAI21X2 U662 ( .A(n601), .B(n603), .C(n835), .Z(n602) );
  HS65_LL_OAI21X2 U663 ( .A(n749), .B(n618), .C(n744), .Z(n617) );
  HS65_LL_IVX4 U664 ( .A(n797), .Z(n936) );
  HS65_LL_IVX4 U665 ( .A(n713), .Z(n714) );
  HS65_LL_IVX4 U666 ( .A(n709), .Z(n710) );
  HS65_LL_OAI21X5 U667 ( .A(N400), .B(n858), .C(n646), .Z(n709) );
  HS65_LL_IVX4 U668 ( .A(n648), .Z(n693) );
  HS65_LL_NAND2X4 U669 ( .A(n805), .B(n893), .Z(n940) );
  HS65_LL_NAND2X7 U670 ( .A(n859), .B(N411), .Z(n534) );
  HS65_LL_NAND2X7 U671 ( .A(N400), .B(n858), .Z(n646) );
  HS65_LL_NAND2X7 U672 ( .A(N523), .B(n836), .Z(n599) );
  HS65_LL_OAI12X2 U673 ( .A(n803), .B(n802), .C(n801), .Z(n921) );
  HS65_LL_NAND2X4 U674 ( .A(N1144), .B(n841), .Z(n833) );
  HS65_LL_OAI12X2 U675 ( .A(n652), .B(n651), .C(n650), .Z(n927) );
  HS65_LL_OAI12X2 U676 ( .A(N523), .B(n700), .C(n699), .Z(n816) );
  HS65_LL_AND2ABX18 U677 ( .A(n791), .B(n944), .Z(N4740) );
  HS65_LL_AND2ABX18 U678 ( .A(n787), .B(n944), .Z(N4739) );
  HS65_LL_AND2ABX18 U679 ( .A(n789), .B(n944), .Z(N4738) );
  HS65_LL_NOR2X5 U680 ( .A(N610), .B(n667), .Z(n972) );
  HS65_LL_NOR2X6 U681 ( .A(n888), .B(N619), .Z(n806) );
  HS65_LL_IVX4 U682 ( .A(N596), .Z(n800) );
  HS65_LL_IVX4 U683 ( .A(N580), .Z(n979) );
  HS65_LL_BFX18 U684 ( .A(N293), .Z(N816) );
  HS65_LL_BFX13 U685 ( .A(N592), .Z(N1066) );
  HS65_LL_NOR2X5 U686 ( .A(N616), .B(N613), .Z(n968) );
  HS65_LL_IVX4 U687 ( .A(N468), .Z(n742) );
  HS65_LL_IVX4 U688 ( .A(N374), .Z(n658) );
  HS65_LL_IVX4 U689 ( .A(N607), .Z(n667) );
  HS65_LL_IVX13 U690 ( .A(N332), .Z(n842) );
  HS65_LL_IVX4 U691 ( .A(N595), .Z(n798) );
  HS65_LL_NOR2X5 U692 ( .A(N610), .B(N607), .Z(n973) );
  HS65_LL_BFX13 U693 ( .A(N549), .Z(N2387) );
  HS65_LL_OAI212X5 U694 ( .A(N574), .B(n644), .C(n664), .D(n643), .E(N2139), 
        .Z(n645) );
  HS65_LL_IVX7 U695 ( .A(n642), .Z(n517) );
  HS65_LL_IVX13 U696 ( .A(n753), .Z(N7604) );
  HS65_LL_IVX13 U697 ( .A(n881), .Z(N8075) );
  HS65_LL_IVX13 U698 ( .A(n759), .Z(N7600) );
  HS65_LL_AOI21X2 U699 ( .A(N625), .B(N118), .C(n889), .Z(n890) );
  HS65_LL_NAND2X7 U700 ( .A(n585), .B(n530), .Z(n975) );
  HS65_LL_AOI21X2 U701 ( .A(n888), .B(n887), .C(n886), .Z(n889) );
  HS65_LL_OA12X4 U702 ( .A(n882), .B(n880), .C(n879), .Z(n881) );
  HS65_LL_AOI12X23 U703 ( .A(N631), .B(N135), .C(n900), .Z(N7626) );
  HS65_LL_IVX13 U704 ( .A(n698), .Z(N7470) );
  HS65_LL_OAI12X3 U705 ( .A(N599), .B(n899), .C(n898), .Z(n900) );
  HS65_LL_MX41X14 U706 ( .D0(n902), .S0(n959), .D1(n901), .S1(n958), .D2(n957), 
        .S2(N173), .D3(n956), .S3(N203), .Z(N7758) );
  HS65_LL_IVX7 U707 ( .A(n960), .Z(n976) );
  HS65_LL_OAI222X5 U708 ( .A(n731), .B(N7432), .C(n897), .D(n734), .E(n882), 
        .F(n894), .Z(n969) );
  HS65_LLS_XOR2X6 U709 ( .A(n555), .B(n554), .Z(n573) );
  HS65_LL_IVX13 U710 ( .A(n719), .Z(N7471) );
  HS65_LL_NAND3X5 U711 ( .A(n762), .B(n761), .C(n760), .Z(n902) );
  HS65_LL_OAI22X4 U712 ( .A(n829), .B(n731), .C(n818), .D(n882), .Z(n689) );
  HS65_LL_AO12X4 U713 ( .A(n806), .B(N122), .C(n697), .Z(n698) );
  HS65_LL_MUX21I1X3 U714 ( .D0(n610), .D1(n609), .S0(n608), .Z(n629) );
  HS65_LLS_XNOR2X3 U715 ( .A(n653), .B(n795), .Z(n915) );
  HS65_LL_OAI12X3 U716 ( .A(n737), .B(n795), .C(n736), .Z(n738) );
  HS65_LL_OAI12X3 U717 ( .A(n677), .B(n795), .C(n676), .Z(n678) );
  HS65_LL_MUXI21X2 U718 ( .D0(n569), .D1(n568), .S0(n567), .Z(n570) );
  HS65_LL_OAI12X3 U719 ( .A(n795), .B(n935), .C(n794), .Z(n796) );
  HS65_LLS_XNOR2X3 U720 ( .A(n627), .B(n626), .Z(n628) );
  HS65_LL_AO12X4 U721 ( .A(n806), .B(N128), .C(n649), .Z(n719) );
  HS65_LL_AOI12X4 U722 ( .A(n745), .B(n943), .C(n941), .Z(n804) );
  HS65_LL_MUXI21X2 U723 ( .D0(n625), .D1(n624), .S0(n623), .Z(n626) );
  HS65_LLS_XNOR2X3 U724 ( .A(n672), .B(n745), .Z(n824) );
  HS65_LL_OAI21X2 U725 ( .A(n592), .B(n595), .C(n591), .Z(n593) );
  HS65_LL_IVX4 U726 ( .A(n543), .Z(n544) );
  HS65_LL_AOI12X23 U727 ( .A(n806), .B(N129), .C(n725), .Z(N7363) );
  HS65_LL_NAND2AX4 U728 ( .A(n548), .B(n693), .Z(n565) );
  HS65_LL_NOR2X5 U729 ( .A(n682), .B(n681), .Z(n712) );
  HS65_LL_AOI21X2 U730 ( .A(n730), .B(n660), .C(n707), .Z(n543) );
  HS65_LL_NOR2X5 U731 ( .A(n537), .B(n538), .Z(n545) );
  HS65_LLS_XNOR2X3 U732 ( .A(n619), .B(n852), .Z(n624) );
  HS65_LL_IVX4 U733 ( .A(n622), .Z(n596) );
  HS65_LL_OAI21X2 U734 ( .A(n835), .B(n603), .C(n602), .Z(n604) );
  HS65_LL_OAI21X2 U735 ( .A(n744), .B(n618), .C(n617), .Z(n619) );
  HS65_LL_AOI12X4 U736 ( .A(n590), .B(n589), .C(n592), .Z(n622) );
  HS65_LL_OAI12X6 U737 ( .A(n794), .B(n936), .C(n561), .Z(n950) );
  HS65_LL_IVX7 U738 ( .A(n729), .Z(n730) );
  HS65_LL_NAND2X5 U739 ( .A(n726), .B(n729), .Z(n536) );
  HS65_LL_OAI12X3 U740 ( .A(n943), .B(n941), .C(n805), .Z(n613) );
  HS65_LLS_XNOR2X3 U741 ( .A(n703), .B(n714), .Z(n595) );
  HS65_LL_OAI12X3 U742 ( .A(n621), .B(n822), .C(n600), .Z(n589) );
  HS65_LL_IVX13 U743 ( .A(n525), .Z(N6716) );
  HS65_LL_OAI12X3 U744 ( .A(n748), .B(n615), .C(n616), .Z(n941) );
  HS65_LL_NOR2X5 U745 ( .A(n542), .B(n541), .Z(n729) );
  HS65_LL_NOR2X5 U746 ( .A(n748), .B(n672), .Z(n943) );
  HS65_LL_NAND2X11 U747 ( .A(n587), .B(n600), .Z(n822) );
  HS65_LL_OAI12X3 U748 ( .A(n599), .B(n713), .C(n684), .Z(n592) );
  HS65_LL_NOR2X5 U749 ( .A(n559), .B(n557), .Z(n739) );
  HS65_LLS_XNOR3X2 U750 ( .A(n582), .B(n581), .C(n580), .Z(n518) );
  HS65_LL_OAI12X3 U751 ( .A(n600), .B(n702), .C(n599), .Z(n603) );
  HS65_LL_OAI12X3 U752 ( .A(n805), .B(n893), .C(n940), .Z(n852) );
  HS65_LL_IVX7 U753 ( .A(n736), .Z(n562) );
  HS65_LL_NAND2X5 U754 ( .A(n616), .B(n612), .Z(n748) );
  HS65_LL_NAND2X5 U755 ( .A(N534), .B(n840), .Z(n600) );
  HS65_LL_NAND2X5 U756 ( .A(n868), .B(N457), .Z(n561) );
  HS65_LL_IVX7 U757 ( .A(n534), .Z(n542) );
  HS65_LL_NOR3X1 U758 ( .A(n922), .B(n921), .C(n920), .Z(n923) );
  HS65_LL_OAI12X3 U759 ( .A(n648), .B(n646), .C(n532), .Z(n691) );
  HS65_LL_OAI21X9 U760 ( .A(N523), .B(n836), .C(n599), .Z(n702) );
  HS65_LL_NOR3X1 U761 ( .A(n811), .B(n810), .C(n809), .Z(n812) );
  HS65_LL_NOR2X5 U762 ( .A(n862), .B(n742), .Z(n559) );
  HS65_LL_IVX7 U763 ( .A(n839), .Z(n840) );
  HS65_LL_NOR2X5 U764 ( .A(n871), .B(n658), .Z(n726) );
  HS65_LL_OAI21X2 U765 ( .A(n659), .B(n658), .C(n657), .Z(n920) );
  HS65_LL_NOR2X5 U766 ( .A(N411), .B(n859), .Z(n541) );
  HS65_LL_NOR2X5 U767 ( .A(N54), .B(n835), .Z(n723) );
  HS65_LL_OAI21X2 U768 ( .A(N323), .B(N372), .C(n841), .Z(n846) );
  HS65_LL_IVX7 U769 ( .A(n835), .Z(n621) );
  HS65_LL_MUXI21X5 U770 ( .D0(N288), .D1(N281), .S0(n853), .Z(n871) );
  HS65_LL_MUX21X4 U771 ( .D0(N264), .D1(N257), .S0(n853), .Z(n531) );
  HS65_LL_MUXI21X2 U772 ( .D0(N217), .D1(N210), .S0(n853), .Z(n869) );
  HS65_LL_IVX7 U773 ( .A(n842), .Z(n841) );
  HS65_LL_OAI12X3 U774 ( .A(n842), .B(N338), .C(N514), .Z(n684) );
  HS65_LL_IVX4 U775 ( .A(N709), .Z(n944) );
  HS65_LL_IVX9 U776 ( .A(n731), .Z(n516) );
  HS65_LL_IVX4 U777 ( .A(N619), .Z(n886) );
  HS65_LL_IVX7 U778 ( .A(N341), .Z(n780) );
  HS65_LL_IVX13 U779 ( .A(N366), .Z(N1139) );
  HS65_LL_IVX13 U780 ( .A(N562), .Z(N1154) );
  HS65_LL_IVX13 U781 ( .A(N338), .Z(N1144) );
  HS65_LL_IVX13 U782 ( .A(N559), .Z(N1155) );
  HS65_LL_IVX13 U783 ( .A(N245), .Z(N1152) );
  HS65_LL_BFX27 U784 ( .A(N299), .Z(N2527) );
  HS65_LL_IVX27 U785 ( .A(N335), .Z(n853) );
  HS65_LL_IVX13 U786 ( .A(N552), .Z(N1153) );
  HS65_LL_IVX13 U787 ( .A(N348), .Z(N1138) );
  HS65_LL_MUX21X18 U788 ( .D0(n892), .D1(n893), .S0(n907), .Z(N7432) );
  HS65_LL_AO222X4 U789 ( .A(n919), .B(n516), .C(n806), .D(N115), .E(n922), .F(
        n885), .Z(n519) );
  HS65_LL_MUX21X9 U790 ( .D0(n976), .D1(n975), .S0(N577), .Z(n980) );
  HS65_LLS_XNOR2X6 U791 ( .A(n571), .B(n570), .Z(n572) );
  HS65_LL_OA12X9 U792 ( .A(n936), .B(n935), .C(n676), .Z(n677) );
  HS65_LL_IVX9 U793 ( .A(n882), .Z(n885) );
  HS65_LL_NAND2AX4 U794 ( .A(n535), .B(n646), .Z(n538) );
  HS65_LL_IVX2 U795 ( .A(n687), .Z(n686) );
  HS65_LL_NAND2AX4 U796 ( .A(n805), .B(n616), .Z(n618) );
  HS65_LLS_XOR3X2 U797 ( .A(n539), .B(n706), .C(n543), .Z(n540) );
  HS65_LL_IVX2 U798 ( .A(N457), .Z(n802) );
  HS65_LL_IVX2 U799 ( .A(N422), .Z(n651) );
  HS65_LL_IVX2 U800 ( .A(n702), .Z(n703) );
  HS65_LL_NOR2X2 U801 ( .A(n680), .B(n722), .Z(n701) );
  HS65_LL_IVX2 U802 ( .A(n748), .Z(n749) );
  HS65_LL_CBI4I1X3 U803 ( .A(n707), .B(N4), .C(n706), .D(n710), .Z(n690) );
  HS65_LL_IVX2 U804 ( .A(N218), .Z(n772) );
  HS65_LL_IVX2 U805 ( .A(N226), .Z(n774) );
  HS65_LL_IVX2 U806 ( .A(N210), .Z(n799) );
  HS65_LL_IVX2 U807 ( .A(N369), .Z(n843) );
  HS65_LL_IVX2 U808 ( .A(N316), .Z(n844) );
  HS65_LL_OAI212X3 U809 ( .A(N265), .B(N597), .C(n771), .D(N598), .E(N400), 
        .Z(n704) );
  HS65_LL_OAI212X3 U810 ( .A(N281), .B(n800), .C(n656), .D(n798), .E(n658), 
        .Z(n657) );
  HS65_LL_IVX2 U811 ( .A(N281), .Z(n656) );
  HS65_LL_IVX2 U812 ( .A(N577), .Z(n977) );
  HS65_LL_IVX2 U813 ( .A(N574), .Z(n664) );
  HS65_LL_NAND2X2 U814 ( .A(n927), .B(n885), .Z(n762) );
  HS65_LL_NAND2X2 U815 ( .A(N113), .B(n806), .Z(n761) );
  HS65_LL_NAND2X2 U816 ( .A(N112), .B(n806), .Z(n674) );
  HS65_LL_NAND2X2 U817 ( .A(n885), .B(n813), .Z(n675) );
  HS65_LL_IVX2 U818 ( .A(N603), .Z(n896) );
  HS65_LL_IVX2 U819 ( .A(N123), .Z(n897) );
  HS65_LL_IVX2 U820 ( .A(n824), .Z(n827) );
  HS65_LL_AOI12X2 U821 ( .A(n707), .B(N4), .C(n706), .Z(n708) );
  HS65_LL_MUX21I1X3 U822 ( .D0(N4), .D1(N4), .S0(n660), .Z(n909) );
  HS65_LL_MUX21I1X3 U823 ( .D0(n695), .D1(n695), .S0(n694), .Z(n912) );
  HS65_LL_AOI12X2 U824 ( .A(n693), .B(n692), .C(n691), .Z(n694) );
  HS65_LL_IVX2 U825 ( .A(n690), .Z(n692) );
  HS65_LL_AOI212X2 U826 ( .A(N257), .B(N289), .C(n855), .D(n854), .E(N335), 
        .Z(n856) );
  HS65_LL_MUX21X4 U827 ( .D0(n687), .D1(n686), .S0(n685), .Z(n829) );
  HS65_LL_NOR2X2 U828 ( .A(n712), .B(n713), .Z(n683) );
  HS65_LL_IVX2 U829 ( .A(n893), .Z(n892) );
  HS65_LL_MUXI21X2 U830 ( .D0(N2527), .D1(N816), .S0(n842), .Z(n893) );
  HS65_LL_IVX2 U831 ( .A(N131), .Z(n655) );
  HS65_LL_IVX2 U832 ( .A(n810), .Z(n654) );
  HS65_LL_IVX2 U833 ( .A(N257), .Z(n855) );
  HS65_LL_IVX2 U834 ( .A(N289), .Z(n854) );
  HS65_LL_OAI212X3 U835 ( .A(N341), .B(N597), .C(n780), .D(N598), .E(N523), 
        .Z(n699) );
  HS65_LL_IVX2 U836 ( .A(N588), .Z(n947) );
  HS65_LL_NAND3X2 U837 ( .A(n548), .B(n545), .C(n544), .Z(n546) );
  HS65_LL_OR2X4 U838 ( .A(n545), .B(n544), .Z(n547) );
  HS65_LL_MUXI41X2 U839 ( .D0(N242), .D1(n631), .D2(N254), .D3(n630), .S0(N400), .S1(n771), .Z(n576) );
  HS65_LL_IVX2 U840 ( .A(n595), .Z(n597) );
  HS65_LL_IVX2 U841 ( .A(N583), .Z(n608) );
  HS65_LL_IVX2 U842 ( .A(n600), .Z(n680) );
  HS65_LL_IVX2 U843 ( .A(n938), .Z(n671) );
  HS65_LL_NOR2X2 U844 ( .A(N457), .B(n868), .Z(n560) );
  HS65_LL_NOR2X2 U845 ( .A(N468), .B(n863), .Z(n557) );
  HS65_LL_IVX2 U846 ( .A(n599), .Z(n682) );
  HS65_LL_NOR2X2 U847 ( .A(n822), .B(n702), .Z(n601) );
  HS65_LL_NAND2AX4 U848 ( .A(N479), .B(n849), .Z(n612) );
  HS65_LL_NAND2X2 U849 ( .A(n710), .B(n707), .Z(n548) );
  HS65_LL_IVX2 U850 ( .A(n615), .Z(n744) );
  HS65_LL_OR2X4 U851 ( .A(N490), .B(n611), .Z(n746) );
  HS65_LL_NAND2AX4 U852 ( .A(n726), .B(n514), .Z(n660) );
  HS65_LL_NAND2X2 U853 ( .A(N389), .B(n531), .Z(n532) );
  HS65_LL_IVX2 U854 ( .A(n950), .Z(n676) );
  HS65_LL_NOR2X2 U855 ( .A(N422), .B(n866), .Z(n737) );
  HS65_LL_NAND2X2 U856 ( .A(n866), .B(N422), .Z(n736) );
  HS65_LL_MUXI21X2 U857 ( .D0(N225), .D1(N218), .S0(n853), .Z(n862) );
  HS65_LL_IVX2 U858 ( .A(n865), .Z(n866) );
  HS65_LL_IVX2 U859 ( .A(n862), .Z(n863) );
  HS65_LL_NAND2X2 U860 ( .A(n871), .B(n658), .Z(n727) );
  HS65_LL_NAND2AX4 U861 ( .A(n849), .B(N479), .Z(n616) );
  HS65_LL_NOR2X2 U862 ( .A(n702), .B(n713), .Z(n590) );
  HS65_LL_NOR2X2 U863 ( .A(n648), .B(n709), .Z(n533) );
  HS65_LL_AND2X4 U864 ( .A(n714), .B(n601), .Z(n620) );
  HS65_LL_IVX2 U865 ( .A(n951), .Z(n934) );
  HS65_LL_OAI212X3 U866 ( .A(N218), .B(n800), .C(n772), .D(n798), .E(n742), 
        .Z(n741) );
  HS65_LL_OAI212X3 U867 ( .A(N226), .B(n800), .C(n774), .D(n798), .E(n651), 
        .Z(n650) );
  HS65_LL_IVX2 U868 ( .A(n679), .Z(n922) );
  HS65_LL_OAI212X3 U869 ( .A(N210), .B(n800), .C(n799), .D(n798), .E(n802), 
        .Z(n801) );
  HS65_LL_NAND2X2 U870 ( .A(n888), .B(n877), .Z(n878) );
  HS65_LL_AO222X4 U871 ( .A(n825), .B(n516), .C(n806), .D(N116), .E(n814), .F(
        n885), .Z(n528) );
  HS65_LL_NAND2X2 U872 ( .A(n646), .B(n690), .Z(n647) );
  HS65_LL_MUXI21X2 U873 ( .D0(n936), .D1(n797), .S0(n796), .Z(n918) );
  HS65_LL_MUXI21X2 U874 ( .D0(n934), .D1(n951), .S0(n678), .Z(n919) );
  HS65_LL_IVX2 U875 ( .A(n739), .Z(n740) );
  HS65_LL_OAI22X1 U876 ( .A(n912), .B(n731), .C(n926), .D(n882), .Z(n697) );
  HS65_LL_PAOI2X3 U877 ( .A(n834), .B(n622), .P(n688), .Z(n942) );
  HS65_LL_IVX2 U878 ( .A(N265), .Z(n771) );
  HS65_LL_IVX2 U879 ( .A(N361), .Z(n781) );
  HS65_LL_NAND3X2 U880 ( .A(n687), .B(n621), .C(n620), .Z(n938) );
  HS65_LL_IVX2 U881 ( .A(n670), .Z(n813) );
  HS65_LL_IVX2 U882 ( .A(n750), .Z(n814) );
  HS65_LL_MX41X4 U883 ( .D0(n902), .S0(n964), .D1(n901), .S1(n963), .D2(n962), 
        .S2(N173), .D3(n961), .S3(N203), .Z(n763) );
  HS65_LL_AOI22X1 U884 ( .A(N40), .B(n966), .C(N91), .D(n965), .Z(n905) );
  HS65_LL_OAI212X3 U885 ( .A(N603), .B(n897), .C(n896), .D(N7432), .E(N599), 
        .Z(n898) );
  HS65_LL_IVX2 U886 ( .A(n820), .Z(n831) );
  HS65_LL_CBI4I6X2 U887 ( .A(N264), .B(N292), .C(n857), .D(n856), .Z(n874) );
  HS65_LL_CBI4I1X3 U888 ( .A(N372), .B(N323), .C(n846), .D(n845), .Z(n847) );
  HS65_LL_IVX2 U889 ( .A(N126), .Z(n733) );
  HS65_LL_AO112X4 U890 ( .A(n723), .B(n822), .C(n722), .D(n731), .Z(n724) );
  HS65_LL_IVX2 U891 ( .A(N34), .Z(n945) );
  HS65_LL_IVX2 U892 ( .A(N88), .Z(n946) );
  HS65_LLS_XNOR3X2 U893 ( .A(n584), .B(n583), .C(n518), .Z(n883) );
  HS65_LL_MX41X14 U894 ( .D0(n520), .S0(n964), .D1(n528), .S1(n963), .D2(n962), 
        .S2(N167), .D3(n961), .S3(N197), .Z(N7755) );
  HS65_LL_OAI212X3 U895 ( .A(N316), .B(N369), .C(n844), .D(n843), .E(n842), 
        .Z(n845) );
  HS65_LL_AO222X4 U896 ( .A(n916), .B(n516), .C(n806), .D(N53), .E(n928), .F(
        n885), .Z(n520) );
  HS65_LL_MX41X14 U897 ( .D0(n969), .S0(n973), .D1(n519), .S1(n974), .D2(n971), 
        .S2(N106), .D3(n972), .S3(N109), .Z(N7736) );
  HS65_LL_AND2X4 U898 ( .A(n924), .B(n923), .Z(n521) );
  HS65_LL_AO222X4 U899 ( .A(n930), .B(n885), .C(n806), .D(N127), .E(n516), .F(
        n910), .Z(n523) );
  HS65_LL_AO222X4 U900 ( .A(n816), .B(n885), .C(n806), .D(N119), .E(n516), .F(
        n821), .Z(n524) );
  HS65_LLS_XNOR3X2 U901 ( .A(N302), .B(N816), .C(n786), .Z(n525) );
  HS65_LL_AND2X4 U902 ( .A(n932), .B(n931), .Z(n527) );
  HS65_LL_MX41X14 U903 ( .D0(n969), .S0(n968), .D1(n519), .S1(n967), .D2(n966), 
        .S2(N106), .D3(n965), .S3(N109), .Z(N7735) );
  HS65_LL_AND2X4 U904 ( .A(n716), .B(n715), .Z(n529) );
  HS65_LL_NAND2X2 U905 ( .A(n885), .B(n883), .Z(n530) );
  HS65_LL_MUXI21X2 U906 ( .D0(N241), .D1(N234), .S0(n853), .Z(n861) );
  HS65_LL_MUXI21X2 U907 ( .D0(n696), .D1(N435), .S0(n861), .Z(n695) );
  HS65_LL_MUX21I1X6 U908 ( .D0(N389), .D1(N389), .S0(n531), .Z(n648) );
  HS65_LL_MUX21X9 U909 ( .D0(N272), .D1(N265), .S0(n853), .Z(n858) );
  HS65_LLS_XOR3X2 U910 ( .A(n695), .B(n693), .C(n709), .Z(n555) );
  HS65_LL_MUX21X9 U911 ( .D0(N280), .D1(N273), .S0(n853), .Z(n859) );
  HS65_LL_NOR2X2 U912 ( .A(n709), .B(n534), .Z(n535) );
  HS65_LL_NOR2X2 U913 ( .A(n709), .B(n536), .Z(n537) );
  HS65_LL_MUXI21X2 U914 ( .D0(n538), .D1(n545), .S0(n726), .Z(n539) );
  HS65_LL_MUXI21X2 U915 ( .D0(n542), .D1(n541), .S0(n514), .Z(n551) );
  HS65_LL_NAND2X2 U916 ( .A(n566), .B(n565), .Z(n549) );
  HS65_LL_NOR2AX3 U917 ( .A(n561), .B(n560), .Z(n797) );
  HS65_LL_MUXI21X2 U918 ( .D0(N209), .D1(N206), .S0(n853), .Z(n954) );
  HS65_LL_MUXI21X2 U919 ( .D0(N446), .D1(n953), .S0(n954), .Z(n951) );
  HS65_LLS_XOR3X2 U920 ( .A(n936), .B(n556), .C(n951), .Z(n571) );
  HS65_LL_MUXI21X2 U921 ( .D0(n557), .D1(n559), .S0(n737), .Z(n558) );
  HS65_LL_MUXI21X2 U922 ( .D0(n950), .D1(n560), .S0(n559), .Z(n564) );
  HS65_LL_MUXI21X2 U923 ( .D0(n950), .D1(n561), .S0(n794), .Z(n563) );
  HS65_LL_MUXI21X2 U924 ( .D0(n564), .D1(n563), .S0(n562), .Z(n568) );
  HS65_LLS_XNOR2X6 U925 ( .A(n573), .B(n572), .Z(n887) );
  HS65_LL_AND2X4 U926 ( .A(N625), .B(N97), .Z(n574) );
  HS65_LL_IVX9 U927 ( .A(N251), .Z(n630) );
  HS65_LL_IVX9 U928 ( .A(N248), .Z(n631) );
  HS65_LL_MUXI41X2 U929 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n651), .S1(N226), .Z(n584) );
  HS65_LL_MUXI41X2 U930 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n658), .S1(N281), .Z(n583) );
  HS65_LL_MUXI41X2 U931 ( .D0(N254), .D1(n630), .D2(N242), .D3(n631), .S0(N411), .S1(N273), .Z(n582) );
  HS65_LL_MUXI41X2 U932 ( .D0(N242), .D1(n631), .D2(N254), .D3(n630), .S0(N389), .S1(n855), .Z(n581) );
  HS65_LL_MUXI41X2 U933 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n696), .S1(N234), .Z(n579) );
  HS65_LL_MUXI41X2 U934 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n742), .S1(N218), .Z(n578) );
  HS65_LL_MUXI41X2 U935 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n802), .S1(N210), .Z(n575) );
  HS65_LLS_XOR3X2 U936 ( .A(n576), .B(n679), .C(n575), .Z(n577) );
  HS65_LLS_XOR3X2 U937 ( .A(n579), .B(n578), .C(n577), .Z(n580) );
  HS65_LL_NAND2AX7 U938 ( .A(N534), .B(n839), .Z(n587) );
  HS65_LL_MUXI21X2 U939 ( .D0(N1139), .D1(n781), .S0(n842), .Z(n835) );
  HS65_LL_MUXI21X5 U940 ( .D0(N1138), .D1(n780), .S0(n842), .Z(n836) );
  HS65_LL_IVX2 U941 ( .A(n836), .Z(n837) );
  HS65_LL_AOI12X2 U942 ( .A(n837), .B(n587), .C(n682), .Z(n586) );
  HS65_LL_AOI12X2 U943 ( .A(n587), .B(N523), .C(n586), .Z(n588) );
  HS65_LLS_XOR3X2 U944 ( .A(n822), .B(n835), .C(n588), .Z(n594) );
  HS65_LL_MUXI21X2 U945 ( .D0(N324), .D1(N331), .S0(n841), .Z(n834) );
  HS65_LL_MUXI21X2 U946 ( .D0(N503), .D1(n688), .S0(n834), .Z(n687) );
  HS65_LL_AOI12X2 U947 ( .A(n596), .B(n595), .C(n620), .Z(n591) );
  HS65_LLS_XOR3X2 U948 ( .A(n594), .B(n686), .C(n593), .Z(n610) );
  HS65_LL_AOI12X2 U949 ( .A(n839), .B(n621), .C(n680), .Z(n598) );
  HS65_LL_AOI12X2 U950 ( .A(n621), .B(N534), .C(n598), .Z(n605) );
  HS65_LLS_XOR3X2 U951 ( .A(n605), .B(n686), .C(n604), .Z(n606) );
  HS65_LL_MUXI21X2 U952 ( .D0(N315), .D1(N308), .S0(n842), .Z(n849) );
  HS65_LL_MUX21X4 U953 ( .D0(N323), .D1(N316), .S0(n842), .Z(n611) );
  HS65_LL_MUX21X4 U954 ( .D0(n616), .D1(n612), .S0(n746), .Z(n614) );
  HS65_LL_MUXI21X2 U955 ( .D0(N302), .D1(N307), .S0(n841), .Z(n805) );
  HS65_LLS_XNOR3X2 U956 ( .A(n614), .B(n892), .C(n613), .Z(n625) );
  HS65_LLS_XNOR2X6 U957 ( .A(n629), .B(n628), .Z(n877) );
  HS65_LL_NAND2X2 U958 ( .A(N625), .B(N94), .Z(n640) );
  HS65_LL_MUXI41X2 U959 ( .D0(N242), .D1(n631), .D2(N254), .D3(n630), .S0(N490), .S1(n844), .Z(n670) );
  HS65_LL_MUXI41X2 U960 ( .D0(N254), .D1(n630), .D2(N242), .D3(n631), .S0(N534), .S1(N351), .Z(n638) );
  HS65_LL_MUXI41X2 U961 ( .D0(N242), .D1(n631), .D2(N254), .D3(n630), .S0(N523), .S1(n780), .Z(n636) );
  HS65_LL_MUXI41X2 U962 ( .D0(n630), .D1(N254), .D2(n631), .D3(N242), .S0(n688), .S1(N324), .Z(n635) );
  HS65_LL_MUXI41X2 U963 ( .D0(N254), .D1(n630), .D2(N242), .D3(n631), .S0(N479), .S1(N308), .Z(n750) );
  HS65_LL_MUXI21X2 U964 ( .D0(N254), .D1(N242), .S0(N816), .Z(n894) );
  HS65_LL_MUXI21X2 U965 ( .D0(N251), .D1(N248), .S0(N302), .Z(n811) );
  HS65_LL_MUXI21X2 U966 ( .D0(N248), .D1(N251), .S0(n781), .Z(n810) );
  HS65_LL_MUXI21X2 U967 ( .D0(N242), .D1(n631), .S0(N514), .Z(n632) );
  HS65_LLS_XOR3X2 U968 ( .A(n811), .B(n810), .C(n632), .Z(n633) );
  HS65_LLS_XOR3X2 U969 ( .A(n750), .B(n894), .C(n633), .Z(n634) );
  HS65_LLS_XOR3X2 U970 ( .A(n636), .B(n635), .C(n634), .Z(n637) );
  HS65_LLS_XOR3X2 U971 ( .A(n670), .B(n638), .C(n637), .Z(n880) );
  HS65_LL_MUX21X4 U972 ( .D0(N179), .D1(N176), .S0(n663), .Z(n643) );
  HS65_LL_BFX18 U973 ( .A(N137), .Z(N2139) );
  HS65_LL_MUXI21X2 U974 ( .D0(n693), .D1(n648), .S0(n647), .Z(n914) );
  HS65_LL_MUXI41X2 U975 ( .D0(n798), .D1(n800), .D2(N598), .D3(N597), .S0(n855), .S1(N389), .Z(n924) );
  HS65_LL_OAI22X1 U976 ( .A(n914), .B(n731), .C(n924), .D(n882), .Z(n649) );
  HS65_LL_MUXI21X2 U977 ( .D0(N598), .D1(N597), .S0(n774), .Z(n652) );
  HS65_LL_AND3X18 U978 ( .A(n762), .B(n761), .C(n760), .Z(N7707) );
  HS65_LL_MUXI21X2 U979 ( .D0(N598), .D1(N597), .S0(n656), .Z(n659) );
  HS65_LL_AO222X4 U980 ( .A(n920), .B(n885), .C(n806), .D(N117), .E(n516), .F(
        n909), .Z(n832) );
  HS65_LL_NOR2AX3 U981 ( .A(N613), .B(N616), .Z(n967) );
  HS65_LL_AND2X4 U982 ( .A(N613), .B(N616), .Z(n966) );
  HS65_LL_NOR2AX3 U983 ( .A(N616), .B(N613), .Z(n965) );
  HS65_LL_NOR3X4 U984 ( .A(N580), .B(n977), .C(n665), .Z(n959) );
  HS65_LL_NOR3X4 U985 ( .A(N577), .B(N580), .C(n665), .Z(n958) );
  HS65_LL_NOR3X4 U986 ( .A(n665), .B(n977), .C(n979), .Z(n957) );
  HS65_LL_NOR3X4 U987 ( .A(N577), .B(n665), .C(n979), .Z(n956) );
  HS65_LL_NOR3X4 U988 ( .A(N574), .B(n663), .C(n665), .Z(n964) );
  HS65_LL_NOR3X4 U989 ( .A(N571), .B(N574), .C(n665), .Z(n963) );
  HS65_LL_NOR3X4 U990 ( .A(n665), .B(n663), .C(n664), .Z(n962) );
  HS65_LL_NOR3X4 U991 ( .A(N571), .B(n665), .C(n664), .Z(n961) );
  HS65_LL_AND2X4 U992 ( .A(N610), .B(n667), .Z(n974) );
  HS65_LL_NOR2AX3 U993 ( .A(N610), .B(n667), .Z(n971) );
  HS65_LL_IVX13 U994 ( .A(n669), .Z(N7015) );
  HS65_LL_IVX13 U995 ( .A(n901), .Z(N7702) );
  HS65_LL_IVX13 U996 ( .A(n519), .Z(N7704) );
  HS65_LL_MX41X14 U997 ( .D0(n969), .S0(n963), .D1(n519), .S1(n964), .D2(N191), 
        .S2(n961), .D3(N161), .S3(n962), .Z(N7757) );
  HS65_LL_NOR2AX3 U998 ( .A(n684), .B(n683), .Z(n685) );
  HS65_LL_MUXI41X2 U999 ( .D0(N597), .D1(N598), .D2(n800), .D3(n798), .S0(N324), .S1(n688), .Z(n818) );
  HS65_LL_MUXI41X2 U1000 ( .D0(N597), .D1(N598), .D2(n800), .D3(n798), .S0(
        N234), .S1(n696), .Z(n926) );
  HS65_LL_MX41X14 U1001 ( .D0(n767), .S0(n968), .D1(n698), .S1(n967), .D2(n966), .S2(N37), .D3(n965), .S3(N43), .Z(N7519) );
  HS65_LL_MUXI21X2 U1002 ( .D0(n798), .D1(n800), .S0(n780), .Z(n700) );
  HS65_LL_MUXI21X2 U1003 ( .D0(n703), .D1(n702), .S0(n701), .Z(n821) );
  HS65_LL_IVX13 U1004 ( .A(n524), .Z(N7467) );
  HS65_LL_MUXI21X2 U1005 ( .D0(n798), .D1(n800), .S0(n771), .Z(n705) );
  HS65_LL_MUXI21X2 U1006 ( .D0(n710), .D1(n709), .S0(n708), .Z(n910) );
  HS65_LL_IVX13 U1007 ( .A(n523), .Z(N7472) );
  HS65_LL_NAND2X2 U1008 ( .A(n806), .B(N130), .Z(n717) );
  HS65_LL_MUXI21X2 U1009 ( .D0(n714), .D1(n713), .S0(n712), .Z(n820) );
  HS65_LL_NAND2X2 U1010 ( .A(n516), .B(n820), .Z(n716) );
  HS65_LL_MUX21X4 U1011 ( .D0(n798), .D1(N598), .S0(N514), .Z(n809) );
  HS65_LL_NAND2X2 U1012 ( .A(n885), .B(n809), .Z(n715) );
  HS65_LL_IVX13 U1013 ( .A(n718), .Z(N7466) );
  HS65_LL_MUXI41X2 U1014 ( .D0(n800), .D1(n798), .D2(N597), .D3(N598), .S0(
        N351), .S1(N534), .Z(n817) );
  HS65_LL_OAI21X3 U1015 ( .A(n817), .B(n882), .C(n724), .Z(n725) );
  HS65_LL_AOI12X2 U1016 ( .A(N4), .B(n514), .C(n726), .Z(n728) );
  HS65_LL_MUXI21X2 U1017 ( .D0(n730), .D1(n729), .S0(n728), .Z(n911) );
  HS65_LL_MUXI41X2 U1018 ( .D0(n800), .D1(n798), .D2(N597), .D3(N598), .S0(
        N273), .S1(N411), .Z(n925) );
  HS65_LL_OA22X4 U1019 ( .A(n911), .B(n731), .C(n925), .D(n882), .Z(n732) );
  HS65_LL_OA12X18 U1020 ( .A(n734), .B(n733), .C(n732), .Z(N7473) );
  HS65_LL_MUXI21X2 U1021 ( .D0(N598), .D1(N597), .S0(n772), .Z(n743) );
  HS65_LL_IVX13 U1022 ( .A(n520), .Z(N7706) );
  HS65_LL_MUXI21X2 U1023 ( .D0(n749), .D1(n748), .S0(n747), .Z(n825) );
  HS65_LL_MX41X14 U1024 ( .D0(n520), .S0(n959), .D1(n528), .S1(n958), .D2(n957), .S2(N167), .D3(n956), .S3(N197), .Z(N7759) );
  HS65_LL_MX41X7 U1025 ( .D0(n698), .S0(n959), .D1(n767), .S1(n958), .D2(n957), 
        .S2(N170), .D3(n956), .S3(N200), .Z(n752) );
  HS65_LL_IVX9 U1026 ( .A(n752), .Z(n753) );
  HS65_LL_MX41X7 U1027 ( .D0(n698), .S0(n964), .D1(n767), .S1(n963), .D2(n962), 
        .S2(N170), .D3(n961), .S3(N200), .Z(n758) );
  HS65_LL_IVX9 U1028 ( .A(n758), .Z(n759) );
  HS65_LL_IVX2 U1029 ( .A(n763), .Z(n764) );
  HS65_LL_IVX13 U1030 ( .A(n764), .Z(N7754) );
  HS65_LL_MX41X14 U1031 ( .D0(n528), .S0(n973), .D1(n520), .S1(n974), .D2(n971), .S2(N103), .D3(n972), .S3(N100), .Z(N7738) );
  HS65_LL_MX41X14 U1032 ( .D0(n524), .S0(n973), .D1(n523), .S1(n974), .D2(n971), .S2(N17), .D3(n972), .S3(N73), .Z(N7517) );
  HS65_LL_MX41X14 U1033 ( .D0(n767), .S0(n973), .D1(n698), .S1(n974), .D2(n971), .S2(N37), .D3(n972), .S3(N43), .Z(N7515) );
  HS65_LL_MX41X14 U1034 ( .D0(n769), .S0(n973), .D1(n768), .S1(n974), .D2(n971), .S2(N70), .D3(n972), .S3(N67), .Z(N7518) );
  HS65_LL_NAND2X14 U1035 ( .A(N27), .B(N31), .Z(N2623) );
  HS65_LL_IVX2 U1036 ( .A(N2623), .Z(n906) );
  HS65_LL_NAND2X14 U1037 ( .A(n906), .B(N83), .Z(N4279) );
  HS65_LL_NAND2X14 U1038 ( .A(n906), .B(N140), .Z(N2590) );
  HS65_LL_MUXI21X2 U1039 ( .D0(N257), .D1(n855), .S0(n771), .Z(n779) );
  HS65_LL_MUXI21X2 U1040 ( .D0(n854), .D1(N289), .S0(N206), .Z(n778) );
  HS65_LL_MUXI21X2 U1041 ( .D0(n772), .D1(N218), .S0(N234), .Z(n773) );
  HS65_LL_MUXI21X2 U1042 ( .D0(n774), .D1(N226), .S0(n773), .Z(n775) );
  HS65_LL_MUXI21X2 U1043 ( .D0(n799), .D1(N210), .S0(n775), .Z(n776) );
  HS65_LLS_XOR3X2 U1044 ( .A(N273), .B(N281), .C(n776), .Z(n777) );
  HS65_LL_XOR3X18 U1045 ( .A(n779), .B(n778), .C(n777), .Z(N6877) );
  HS65_LL_MUXI21X2 U1046 ( .D0(n780), .D1(N341), .S0(N351), .Z(n785) );
  HS65_LL_MUXI21X2 U1047 ( .D0(n781), .D1(N361), .S0(N324), .Z(n784) );
  HS65_LL_MUXI21X2 U1048 ( .D0(n843), .D1(N369), .S0(N308), .Z(n782) );
  HS65_LL_MUXI21X2 U1049 ( .D0(N316), .D1(n844), .S0(n782), .Z(n783) );
  HS65_LLS_XOR3X2 U1050 ( .A(n785), .B(n784), .C(n783), .Z(n786) );
  HS65_LL_NAND2X14 U1051 ( .A(N556), .B(N386), .Z(N2061) );
  HS65_LL_AOI212X2 U1052 ( .A(N23), .B(N588), .C(N79), .D(n947), .E(N2623), 
        .Z(n787) );
  HS65_LL_BFX27 U1053 ( .A(N141), .Z(N709) );
  HS65_LL_AOI212X2 U1054 ( .A(N81), .B(N588), .C(N26), .D(n947), .E(N2623), 
        .Z(n789) );
  HS65_LL_AOI212X2 U1055 ( .A(N80), .B(N588), .C(N82), .D(n947), .E(N2623), 
        .Z(n791) );
  HS65_LL_AOI212X2 U1056 ( .A(N25), .B(N588), .C(N24), .D(n947), .E(N2623), 
        .Z(n793) );
  HS65_LL_AND2ABX18 U1057 ( .A(n793), .B(n944), .Z(N4737) );
  HS65_LL_MUXI21X2 U1058 ( .D0(N598), .D1(N597), .S0(n799), .Z(n803) );
  HS65_LL_IVX13 U1059 ( .A(n522), .Z(N7705) );
  HS65_LL_IVX13 U1060 ( .A(n807), .Z(N7700) );
  HS65_LL_NAND4ABX3 U1061 ( .A(n814), .B(n813), .C(n894), .D(n812), .Z(n815)
         );
  HS65_LL_IVX13 U1062 ( .A(N358), .Z(N1145) );
  HS65_LL_NOR4ABX2 U1063 ( .A(n823), .B(n893), .C(n822), .D(n821), .Z(n828) );
  HS65_LL_NOR4ABX2 U1064 ( .A(n828), .B(n827), .C(n826), .D(n825), .Z(n830) );
  HS65_LL_AND3X18 U1065 ( .A(n831), .B(n830), .C(n829), .Z(N7504) );
  HS65_LL_IVX13 U1066 ( .A(n832), .Z(N7365) );
  HS65_LL_MX41X14 U1067 ( .D0(n969), .S0(n958), .D1(n519), .S1(n959), .D2(N161), .S2(n957), .D3(n956), .S3(N191), .Z(N7761) );
  HS65_LL_MX41X14 U1068 ( .D0(n719), .S0(n964), .D1(n718), .S1(n963), .D2(n962), .S2(N146), .D3(n961), .S3(N149), .Z(N7603) );
  HS65_LL_MX41X14 U1069 ( .D0(n528), .S0(n968), .D1(n520), .S1(n967), .D2(n966), .S2(N103), .D3(n965), .S3(N100), .Z(N7741) );
  HS65_LL_MX41X14 U1070 ( .D0(n901), .S0(n973), .D1(n902), .S1(n974), .D2(n971), .S2(N40), .D3(n972), .S3(N91), .Z(N7739) );
  HS65_LL_NAND2AX14 U1071 ( .A(N591), .B(N27), .Z(N2060) );
  HS65_LL_MUXI21X2 U1072 ( .D0(N331), .D1(n834), .S0(n833), .Z(n851) );
  HS65_LL_MUXI21X2 U1073 ( .D0(n837), .D1(n836), .S0(n835), .Z(n838) );
  HS65_LL_MUXI21X2 U1074 ( .D0(n840), .D1(n839), .S0(n838), .Z(n848) );
  HS65_LLS_XOR3X2 U1075 ( .A(n849), .B(n848), .C(n847), .Z(n850) );
  HS65_LL_XOR3X18 U1076 ( .A(n852), .B(n851), .C(n850), .Z(N7474) );
  HS65_LL_AOI12X2 U1077 ( .A(N264), .B(N292), .C(n853), .Z(n857) );
  HS65_LL_IVX2 U1078 ( .A(n859), .Z(n860) );
  HS65_LL_MUXI21X2 U1079 ( .D0(n860), .D1(n859), .S0(n858), .Z(n873) );
  HS65_LL_MUXI21X2 U1080 ( .D0(n863), .D1(n862), .S0(n861), .Z(n864) );
  HS65_LL_MUXI21X2 U1081 ( .D0(n866), .D1(n865), .S0(n864), .Z(n867) );
  HS65_LL_MUXI21X2 U1082 ( .D0(n869), .D1(n868), .S0(n867), .Z(n870) );
  HS65_LLS_XOR3X2 U1083 ( .A(n871), .B(n954), .C(n870), .Z(n872) );
  HS65_LL_XOR3X18 U1084 ( .A(n874), .B(n873), .C(n872), .Z(N7476) );
  HS65_LL_AND2ABX18 U1085 ( .A(N1153), .B(N1154), .Z(N1140) );
  HS65_LL_NAND4ABX3 U1086 ( .A(N6716), .B(N2061), .C(N1140), .D(n875), .Z(n876) );
  HS65_LL_AND3ABCX18 U1087 ( .A(N7474), .B(N7476), .C(n876), .Z(N7703) );
  HS65_LL_IVX2 U1088 ( .A(n883), .Z(n884) );
  HS65_LL_NAND2X2 U1089 ( .A(n885), .B(n884), .Z(n891) );
  HS65_LL_NAND2X14 U1090 ( .A(n891), .B(n890), .Z(N8076) );
  HS65_LL_MUXI21X2 U1091 ( .D0(n893), .D1(n892), .S0(N132), .Z(n895) );
  HS65_LL_MUXI21X2 U1092 ( .D0(n895), .D1(n894), .S0(n896), .Z(n899) );
  HS65_LL_NAND2X2 U1093 ( .A(n968), .B(n901), .Z(n904) );
  HS65_LL_NAND2X2 U1094 ( .A(n967), .B(n902), .Z(n903) );
  HS65_LL_OR3ABCX18 U1095 ( .A(n905), .B(n904), .C(n903), .Z(N7742) );
  HS65_LL_MUXI21X20 U1096 ( .D0(n908), .D1(n485), .S0(N132), .Z(N7698) );
  HS65_LL_NOR4ABX2 U1097 ( .A(n912), .B(n911), .C(n910), .D(n909), .Z(n913) );
  HS65_LL_NAND4ABX3 U1098 ( .A(n916), .B(n915), .C(n914), .D(n913), .Z(n917)
         );
  HS65_LL_AND3ABCX18 U1099 ( .A(n919), .B(n918), .C(n917), .Z(N7503) );
  HS65_LL_NAND4ABX3 U1100 ( .A(n928), .B(n927), .C(n926), .D(n925), .Z(n929)
         );
  HS65_LL_IVX2 U1101 ( .A(n929), .Z(n932) );
  HS65_LL_IVX2 U1102 ( .A(n930), .Z(n931) );
  HS65_LL_AND2X27 U1103 ( .A(n937), .B(n949), .Z(N6648) );
  HS65_LL_NOR3AX2 U1104 ( .A(n943), .B(n938), .C(n940), .Z(n939) );
  HS65_LL_BFX27 U1105 ( .A(n939), .Z(N6643) );
  HS65_LL_AO112X27 U1106 ( .A(n943), .B(n942), .C(n941), .D(n940), .Z(N6927)
         );
  HS65_LL_IVX27 U1107 ( .A(N2387), .Z(N1141) );
  HS65_LL_NOR2AX25 U1108 ( .A(N145), .B(n944), .Z(N1147) );
  HS65_LL_AO212X27 U1109 ( .A(n947), .B(n946), .C(N588), .D(n945), .E(N2623), 
        .Z(N4275) );
  HS65_LL_IVX13 U1110 ( .A(N2527), .Z(N3613) );
  HS65_LL_IVX40 U1111 ( .A(N545), .Z(N1137) );
  HS65_LL_BFX62 U1112 ( .A(N1), .Z(N2309) );
  HS65_LL_AND2X18 U1113 ( .A(N2309), .B(N373), .Z(N0) );
  HS65_LL_MX41X14 U1114 ( .D0(n522), .S0(n964), .D1(n807), .S1(n963), .D2(n962), .S2(N164), .D3(n961), .S3(N194), .Z(N7756) );
  HS65_LL_MX41X14 U1115 ( .D0(n522), .S0(n959), .D1(n807), .S1(n958), .D2(n957), .S2(N164), .D3(n956), .S3(N194), .Z(N7760) );
  HS65_LL_MX41X14 U1116 ( .D0(n807), .S0(n968), .D1(n522), .S1(n967), .D2(n966), .S2(N49), .D3(n965), .S3(N46), .Z(N7740) );
  HS65_LL_MX41X14 U1117 ( .D0(n807), .S0(n973), .D1(n522), .S1(n974), .D2(n971), .S2(N49), .D3(n972), .S3(N46), .Z(N7737) );
  HS65_LL_MX41X14 U1118 ( .D0(n517), .S0(n967), .D1(n976), .S1(n968), .D2(N64), 
        .S2(n966), .D3(n965), .S3(N14), .Z(N8124) );
  HS65_LL_MX41X14 U1119 ( .D0(n523), .S0(n964), .D1(n524), .S1(n963), .D2(n962), .S2(N152), .D3(n961), .S3(N155), .Z(N7602) );
  HS65_LL_MX41X14 U1120 ( .D0(n517), .S0(n974), .D1(n976), .S1(n973), .D2(N14), 
        .S2(n972), .D3(N64), .S3(n971), .Z(N8123) );
  HS65_LL_MUX21X4 U1121 ( .D0(N179), .D1(N176), .S0(n977), .Z(n978) );
  HS65_LL_OAI212X20 U1122 ( .A(N580), .B(n980), .C(n979), .D(n978), .E(N2139), 
        .Z(N8128) );
endmodule

